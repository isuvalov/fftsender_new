library	ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

package regs_pack is	

constant FIXPOINT:natural:=5;

type Trx2tx_wires is record
	new_request_received: std_logic;
	number_of_req:std_logic_vector(7 downto 0);
	request_type:std_logic_vector(7 downto 0);
	infinity_measure:std_logic;
	measure_time:std_logic_vector(15 downto 0);  --# in seconds
end record Trx2tx_wires;
							  


end regs_pack;
package body regs_pack is 
	


end package body regs_pack;

