---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
--  version   : $Version: 1.0 $ 
--  revision    : $Revision: 1.1.1.1 $ 
--  designer name   : $Author: jzhang $ 
--  company name    : altera corp.
--  company address : 101 innovation drive
--                      san jose, california 95134
--                      u.s.a.
-- 
--  copyright altera corp. 2003
-- 
-- 
--  $Header: /ipbu/cvs/dsp/projects/FFT/src/rtl/lib/asj_fft_cnt_ctrl.vhd,v 1.1.1.1 2005/12/08 01:14:15 jzhang Exp $ 
--  $log$ 
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all; 
library work;
use work.fft_pack.all;

entity asj_fft_cnt_ctrl is
  generic(
            nps : integer :=256;
            mpr : integer :=16;
            apr : integer :=6;
            abuspr : integer :=24; --4*apr
            rbuspr : integer :=64; --4*mpr
            cbuspr : integer :=128 --2*4*mpr
          );
  port(     clk             : in std_logic;
            sel_anb_in      : in std_logic;
            sel_anb_ram     : in std_logic;
            sel_anb_addr    : in std_logic;
            data_rdy        : in std_logic;
            wraddr_i0_sw    : in std_logic_vector(apr-1 downto 0);
            wraddr_i1_sw    : in std_logic_vector(apr-1 downto 0);
            wraddr_i2_sw    : in std_logic_vector(apr-1 downto 0);
            wraddr_i3_sw    : in std_logic_vector(apr-1 downto 0);
            wraddr0_sw    : in std_logic_vector(apr-1 downto 0);
            wraddr1_sw    : in std_logic_vector(apr-1 downto 0);
            wraddr2_sw    : in std_logic_vector(apr-1 downto 0);
            wraddr3_sw    : in std_logic_vector(apr-1 downto 0);
            rdaddr0_sw    : in std_logic_vector(apr-1 downto 0);
            rdaddr1_sw    : in std_logic_vector(apr-1 downto 0);
            rdaddr2_sw    : in std_logic_vector(apr-1 downto 0);
            rdaddr3_sw    : in std_logic_vector(apr-1 downto 0);
            ram_data_in0_sw  : in std_logic_vector(2*mpr-1 downto 0);
            ram_data_in1_sw  : in std_logic_vector(2*mpr-1 downto 0);
            ram_data_in2_sw  : in std_logic_vector(2*mpr-1 downto 0);
            ram_data_in3_sw  : in std_logic_vector(2*mpr-1 downto 0);
            i_ram_data_in0_sw  : in std_logic_vector(2*mpr-1 downto 0);
            i_ram_data_in1_sw  : in std_logic_vector(2*mpr-1 downto 0);
            i_ram_data_in2_sw  : in std_logic_vector(2*mpr-1 downto 0);
            i_ram_data_in3_sw  : in std_logic_vector(2*mpr-1 downto 0);
            a_ram_data_out_bus  : in std_logic_vector(cbuspr-1 downto 0);
            b_ram_data_out_bus  : in std_logic_vector(cbuspr-1 downto 0);
            a_ram_data_in_bus  : out std_logic_vector(cbuspr-1 downto 0);
            b_ram_data_in_bus  : out std_logic_vector(cbuspr-1 downto 0);
            wraddress_a_bus   : out std_logic_vector(abuspr-1 downto 0);
            wraddress_b_bus   : out std_logic_vector(abuspr-1 downto 0);
            rdaddress_a_bus   : out std_logic_vector(abuspr-1 downto 0);
            rdaddress_b_bus   : out std_logic_vector(abuspr-1 downto 0);
            ram_data_out0    : out std_logic_vector(2*mpr-1 downto 0);
            ram_data_out1    : out std_logic_vector(2*mpr-1 downto 0);
            ram_data_out2    : out std_logic_vector(2*mpr-1 downto 0);
            ram_data_out3    : out std_logic_vector(2*mpr-1 downto 0)
            
      );
end asj_fft_cnt_ctrl;

architecture cnt_sw of asj_fft_cnt_ctrl is


begin
  
sel_input_ab : process(clk,sel_anb_in,wraddr_i0_sw,wraddr_i1_sw,wraddr_i2_sw,wraddr_i3_sw,
wraddr0_sw,wraddr1_sw,wraddr2_sw,wraddr3_sw) is
    begin
      if(rising_edge(clk)) then
        if (sel_anb_in='1') then
            wraddress_a_bus <= wraddr_i0_sw & wraddr_i1_sw & wraddr_i2_sw & wraddr_i3_sw;
            wraddress_b_bus <= wraddr0_sw & wraddr1_sw & wraddr2_sw & wraddr3_sw;
        else
            wraddress_b_bus <= wraddr_i0_sw & wraddr_i1_sw & wraddr_i2_sw & wraddr_i3_sw;
            wraddress_a_bus <= wraddr0_sw & wraddr1_sw & wraddr2_sw & wraddr3_sw;
        end if;       
      end if;
    end process sel_input_ab;
    

    
sel_ram_ab : process(clk,sel_anb_in,i_ram_data_in0_sw,ram_data_in0_sw,i_ram_data_in1_sw,ram_data_in1_sw,i_ram_data_in2_sw,ram_data_in2_sw,i_ram_data_in3_sw,ram_data_in3_sw) is
    begin
      if(rising_edge(clk)) then
        if(sel_anb_in='1') then
            a_ram_data_in_bus <= i_ram_data_in0_sw & i_ram_data_in1_sw & i_ram_data_in2_sw & i_ram_data_in3_sw;
            b_ram_data_in_bus <= ram_data_in0_sw & ram_data_in1_sw & ram_data_in2_sw & ram_data_in3_sw;
        else
            b_ram_data_in_bus <= i_ram_data_in0_sw & i_ram_data_in1_sw & i_ram_data_in2_sw & i_ram_data_in3_sw;
            a_ram_data_in_bus <= ram_data_in0_sw & ram_data_in1_sw & ram_data_in2_sw & ram_data_in3_sw;
        end if;       
      end if;
    end process sel_ram_ab;
    
    
sel_ram_data : process(clk,sel_anb_ram,b_ram_data_out_bus,a_ram_data_out_bus) is
    begin
      if(rising_edge(clk)) then
        if(sel_anb_ram='1') then
            ram_data_out0 <= b_ram_data_out_bus(8*mpr-1 downto 6*mpr);
            ram_data_out1 <= b_ram_data_out_bus(6*mpr-1 downto 4*mpr);
            ram_data_out2 <= b_ram_data_out_bus(4*mpr-1 downto 2*mpr);
            ram_data_out3 <= b_ram_data_out_bus(2*mpr-1 downto 0);
        else
            ram_data_out0 <= a_ram_data_out_bus(8*mpr-1 downto 6*mpr);
            ram_data_out1 <= a_ram_data_out_bus(6*mpr-1 downto 4*mpr);
            ram_data_out2 <= a_ram_data_out_bus(4*mpr-1 downto 2*mpr);
            ram_data_out3 <= a_ram_data_out_bus(2*mpr-1 downto 0);
        end if;       
      end if;
    end process sel_ram_data;
    
  sel_ram_addr : process(clk,sel_anb_addr,rdaddr0_sw, rdaddr1_sw ,rdaddr2_sw ,rdaddr3_sw) is
    begin
      if(rising_edge(clk)) then
        if(sel_anb_addr='1') then
            rdaddress_b_bus <= rdaddr0_sw & rdaddr1_sw & rdaddr2_sw & rdaddr3_sw;
            rdaddress_a_bus <= (others=>'0');
        else
            rdaddress_a_bus <= rdaddr0_sw & rdaddr1_sw & rdaddr2_sw & rdaddr3_sw;
            rdaddress_b_bus <= (others=>'0');
        end if;       
      end if;
    end process sel_ram_addr;

  
end cnt_sw;











