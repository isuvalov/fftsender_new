library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;

entity cpp_response2vhdl is
	 port(
		 reset: in std_logic;
		 ce : in std_logic;
		 clk : in std_logic;
		 can_go: in std_logic; --# see falling edge of recieved dv

		 dv_o: out std_logic;
		 data_o: out std_logic_vector(7 downto 0)
	     );
end cpp_response2vhdl;


architecture cpp_response2vhdl of cpp_response2vhdl is

signal delay_cnt:std_logic_vector(3 downto 0):=(others=>'1');
signal cnt:integer:=0;

type Tseq_array0 is array (0 to 42+16-1) of std_logic_vector(7 downto 0);
constant seq_array0:Tseq_array0:=(x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"16", x"ea", x"ca", x"09", x"3a", x"08", x"00", x"45", x"00", x"00", x"1f", x"57", x"ac", x"00", x"00", x"80", x"11", x"21", x"74", x"c0", x"a8", x"01", x"06", x"ff", x"ff", x"ff", x"ff", x"e2", x"ce", x"ec", x"be", x"00", x"0b", x"14", x"9c",
x"A5", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");

type Tseq_array1 is array (0 to 42+5-1) of std_logic_vector(7 downto 0);
constant seq_array1:Tseq_array1:=(x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"16", x"ea", x"ca", x"09", x"3a", x"08", x"00", x"45", x"00", x"00", x"1f", x"57", x"ac", x"00", x"00", x"80", x"11", x"21", x"74", x"c0", x"a8", x"01", x"06", x"ff", x"ff", x"ff", x"ff", x"e2", x"ce", x"ec", x"be", x"00", x"0b", x"14", x"9c",
x"A5", x"02", x"02", x"00", x"04");

type Tseq_array2 is array (0 to 42+10248-1) of std_logic_vector(7 downto 0);
constant seq_array2:Tseq_array2:=(x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"16", x"ea", x"ca", x"09", x"3a", x"08", x"00", x"45", x"00", x"00", x"1f", x"57", x"ac", x"00", x"00", x"80", x"11", x"21", x"74", x"c0", x"a8", x"01", x"06", x"ff", x"ff", x"ff", x"ff", x"e2", x"ce", x"ec", x"be", x"00", x"0b", x"14", x"9c",
x"A5", x"03", x"01", x"00", x"02", x"00", x"5A", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"0A", x"00", x"00", x"00", x"00", x"14", x"00", x"00", x"00", x"00", x"1E", x"00", x"00", x"00", x"00", x"28", x"00", x"00", x"00", x"00", x"32", x"00", x"00", x"00", x"00", x"3C", x"00", x"00", x"00", x"00", x"46", x"00", x"00", x"00", x"00", x"50", x"00", x"00", x"00", x"00", x"5A", x"00", x"00", x"00", x"00", x"64", x"00", x"00", x"00", x"00", x"6E", x"00", x"00", x"00", x"00", x"78", x"00", x"00", x"00", x"00", x"82", x"00", x"00", x"00", x"00", x"8C", x"00", x"00", x"00", x"00", x"96", x"00", x"00", x"00", x"00", x"A0", x"00", x"00", x"00", x"00", x"AA", x"00", x"00", x"00", x"00", x"B4", x"00", x"00", x"00", x"00", x"BE", x"00", x"00", x"00", x"00", x"C8", x"00", x"00", x"00", x"00", x"D2", x"00", x"00", x"00", x"00", x"DC", x"00", x"00", x"00", x"00", x"E6", x"00", x"00", x"00", x"00", x"F0", x"00", x"00", x"00", x"00", x"FA", x"00", x"00", x"00", x"01", x"04", x"00", x"00", x"00", x"01", x"0E", x"00", x"00", x"00", x"01", x"18", x"00", x"00", x"00", x"01", x"22", x"00", x"00", x"00", x"01", x"2C", x"00", x"00", x"00", x"01", x"36", x"00", x"00", x"00", x"01", x"40", x"00", x"00", x"00", x"01", x"4A", x"00", x"00", x"00", x"01", x"54", x"00", x"00", x"00", x"01", x"5E", x"00", x"00", x"00", x"01", x"68", x"00", x"00", x"00", x"01", x"72", x"00", x"00", x"00", x"01", x"7C", x"00", x"00", x"00", x"01", x"86", x"00", x"00", x"00", x"01", x"90", x"00", x"00", x"00", x"01", x"9A", x"00", x"00", x"00", x"01", x"A4", x"00", x"00", x"00", x"01", x"AE", x"00", x"00", x"00", x"01", x"B8", x"00", x"00", x"00", x"01", x"C2", x"00", x"00", x"00", x"01", x"CC", x"00", x"00", x"00", x"01", x"D6", x"00", x"00", x"00", x"01", x"E0", x"00", x"00", x"00", x"01", x"EA", x"00", x"00", x"00", x"01", x"F4", x"00", x"00", x"00", x"01", x"FE", x"00", x"00", x"00", x"02", x"08", x"00", x"00", x"00", x"02", x"12", x"00", x"00", x"00", x"02", x"1C", x"00", x"00", x"00", x"02", x"26", x"00", x"00", x"00", x"02", x"30", x"00", x"00", x"00", x"02", x"3A", x"00", x"00", x"00", x"02", x"44", x"00", x"00", x"00", x"02", x"4E", x"00", x"00", x"00", x"02", x"58", x"00", x"00", x"00", x"02", x"62", x"00", x"00", x"00", x"02", x"6C", x"00", x"00", x"00", x"02", x"76", x"00", x"00", x"00", x"02", x"80", x"00", x"00", x"00", x"02", x"8A", x"00", x"00", x"00", x"02", x"94", x"00", x"00", x"00", x"02", x"9E", x"00", x"00", x"00", x"02", x"A8", x"00", x"00", x"00", x"02", x"B2", x"00", x"00", x"00", x"02", x"BC", x"00", x"00", x"00", x"02", x"C6", x"00", x"00", x"00", x"02", x"D0", x"00", x"00", x"00", x"02", x"DA", x"00", x"00", x"00", x"02", x"E4", x"00", x"00", x"00", x"02", x"EE", x"00", x"00", x"00", x"02", x"F8", x"00", x"00", x"00", x"03", x"02", x"00", x"00", x"00", x"03", x"0C", x"00", x"00", x"00", x"03", x"16", x"00", x"00", x"00", x"03", x"20", x"00", x"00", x"00", x"03", x"2A", x"00", x"00", x"00", x"03", x"34", x"00", x"00", x"00", x"03", x"3E", x"00", x"00", x"00", x"03", x"48", x"00", x"00", x"00", x"03", x"52", x"00", x"00", x"00", x"03", x"5C", x"00", x"00", x"00", x"03", x"66", x"00", x"00", x"00", x"03", x"70", x"00", x"00", x"00", x"03", x"7A", x"00", x"00", x"00", x"03", x"84", x"00", x"00", x"00", x"03", x"8E", x"00", x"00", x"00", x"03", x"98", x"00", x"00", x"00", x"03", x"A2", x"00", x"00", x"00", x"03", x"AC", x"00", x"00", x"00", x"03", x"B6", x"00", x"00", x"00", x"03", x"C0", x"00", x"00", x"00", x"03", x"CA", x"00", x"00", x"00", x"03", x"D4", x"00", x"00", x"00", x"03", x"DE", x"00", x"00", x"00", x"03", x"E8", x"00", x"00", x"00", x"03", x"F2", x"00", x"00", x"00", x"03", x"FC", x"00", x"00", x"00", x"04", x"06", x"00", x"00", x"00", x"04", x"10", x"00", x"00", x"00", x"04", x"1A", x"00", x"00", x"00", x"04", x"24", x"00", x"00", x"00", x"04", x"2E", x"00", x"00", x"00", x"04", x"38", x"00", x"00", x"00", x"04", x"42", x"00", x"00", x"00", x"04", x"4C", x"00", x"00", x"00", x"04", x"56", x"00", x"00", x"00", x"04", x"60", x"00", x"00", x"00", x"04", x"6A", x"00", x"00", x"00", x"04", x"74", x"00", x"00", x"00", x"04", x"7E", x"00", x"00", x"00", x"04", x"88", x"00", x"00", x"00", x"04", x"92", x"00", x"00", x"00", x"04", x"9C", x"00", x"00", x"00", x"04", x"A6", x"00", x"00", x"00", x"04", x"B0", x"00", x"00", x"00", x"04", x"BA", x"00", x"00", x"00", x"04", x"C4", x"00", x"00", x"00", x"04", x"CE", x"00", x"00", x"00", x"04", x"D8", x"00", x"00", x"00", x"04", x"E2", x"00", x"00", x"00", x"04", x"EC", x"00", x"00", x"00", x"04", x"F6", x"00", x"00", x"00", x"05", x"00", x"00", x"00", x"00", x"05", x"0A", x"00", x"00", x"00", x"05", x"14", x"00", x"00", x"00", x"05", x"1E", x"00", x"00", x"00", x"05", x"28", x"00", x"00", x"00", x"05", x"32", x"00", x"00", x"00", x"05", x"3C", x"00", x"00", x"00", x"05", x"46", x"00", x"00", x"00", x"05", x"50", x"00", x"00", x"00", x"05", x"5A", x"00", x"00", x"00", x"05", x"64", x"00", x"00", x"00", x"05", x"6E", x"00", x"00", x"00", x"05", x"78", x"00", x"00", x"00", x"05", x"82", x"00", x"00", x"00", x"05", x"8C", x"00", x"00", x"00", x"05", x"96", x"00", x"00", x"00", x"05", x"A0", x"00", x"00", x"00", x"05", x"AA", x"00", x"00", x"00", x"05", x"B4", x"00", x"00", x"00", x"05", x"BE", x"00", x"00", x"00", x"05", x"C8", x"00", x"00", x"00", x"05", x"D2", x"00", x"00", x"00", x"05", x"DC", x"00", x"00", x"00", x"05", x"E6", x"00", x"00", x"00", x"05", x"F0", x"00", x"00", x"00", x"05", x"FA", x"00", x"00", x"00", x"06", x"04", x"00", x"00", x"00", x"06", x"0E", x"00", x"00", x"00", x"06", x"18", x"00", x"00", x"00", x"06", x"22", x"00", x"00", x"00", x"06", x"2C", x"00", x"00", x"00", x"06", x"36", x"00", x"00", x"00", x"06", x"40", x"00", x"00", x"00", x"06", x"4A", x"00", x"00", x"00", x"06", x"54", x"00", x"00", x"00", x"06", x"5E", x"00", x"00", x"00", x"06", x"68", x"00", x"00", x"00", x"06", x"72", x"00", x"00", x"00", x"06", x"7C", x"00", x"00", x"00", x"06", x"86", x"00", x"00", x"00", x"06", x"90", x"00", x"00", x"00", x"06", x"9A", x"00", x"00", x"00", x"06", x"A4", x"00", x"00", x"00", x"06", x"AE", x"00", x"00", x"00", x"06", x"B8", x"00", x"00", x"00", x"06", x"C2", x"00", x"00", x"00", x"06", x"CC", x"00", x"00", x"00", x"06", x"D6", x"00", x"00", x"00", x"06", x"E0", x"00", x"00", x"00", x"06", x"EA", x"00", x"00", x"00", x"06", x"F4", x"00", x"00", x"00", x"06", x"FE", x"00", x"00", x"00", x"07", x"08", x"00", x"00", x"00", x"07", x"12", x"00", x"00", x"00", x"07", x"1C", x"00", x"00", x"00", x"07", x"26", x"00", x"00", x"00", x"07", x"30", x"00", x"00", x"00", x"07", x"3A", x"00", x"00", x"00", x"07", x"44", x"00", x"00", x"00", x"07", x"4E", x"00", x"00", x"00", x"07", x"58", x"00", x"00", x"00", x"07", x"62", x"00", x"00", x"00", x"07", x"6C", x"00", x"00", x"00", x"07", x"76", x"00", x"00", x"00", x"07", x"80", x"00", x"00", x"00", x"07", x"8A", x"00", x"00", x"00", x"07", x"94", x"00", x"00", x"00", x"07", x"9E", x"00", x"00", x"00", x"07", x"A8", x"00", x"00", x"00", x"07", x"B2", x"00", x"00", x"00", x"07", x"BC", x"00", x"00", x"00", x"07", x"C6", x"00", x"00", x"00", x"07", x"D0", x"00", x"00", x"00", x"07", x"DA", x"00", x"00", x"00", x"07", x"E4", x"00", x"00", x"00", x"07", x"EE", x"00", x"00", x"00", x"07", x"F8", x"00", x"00", x"00", x"08", x"02", x"00", x"00", x"00", x"08", x"0C", x"00", x"00", x"00", x"08", x"16", x"00", x"00", x"00", x"08", x"20", x"00", x"00", x"00", x"08", x"2A", x"00", x"00", x"00", x"08", x"34", x"00", x"00", x"00", x"08", x"3E", x"00", x"00", x"00", x"08", x"48", x"00", x"00", x"00", x"08", x"52", x"00", x"00", x"00", x"08", x"5C", x"00", x"00", x"00", x"08", x"66", x"00", x"00", x"00", x"08", x"70", x"00", x"00", x"00", x"08", x"7A", x"00", x"00", x"00", x"08", x"84", x"00", x"00", x"00", x"08", x"8E", x"00", x"00", x"00", x"08", x"98", x"00", x"00", x"00", x"08", x"A2", x"00", x"00", x"00", x"08", x"AC", x"00", x"00", x"00", x"08", x"B6", x"00", x"00", x"00", x"08", x"C0", x"00", x"00", x"00", x"08", x"CA", x"00", x"00", x"00", x"08", x"D4", x"00", x"00", x"00", x"08", x"DE", x"00", x"00", x"00", x"08", x"E8", x"00", x"00", x"00", x"08", x"F2", x"00", x"00", x"00", x"08", x"FC", x"00", x"00", x"00", x"09", x"06", x"00", x"00", x"00", x"09", x"10", x"00", x"00", x"00", x"09", x"1A", x"00", x"00", x"00", x"09", x"24", x"00", x"00", x"00", x"09", x"2E", x"00", x"00", x"00", x"09", x"38", x"00", x"00", x"00", x"09", x"42", x"00", x"00", x"00", x"09", x"4C", x"00", x"00", x"00", x"09", x"56", x"00", x"00", x"00", x"09", x"60", x"00", x"00", x"00", x"09", x"6A", x"00", x"00", x"00", x"09", x"74", x"00", x"00", x"00", x"09", x"7E", x"00", x"00", x"00", x"09", x"88", x"00", x"00", x"00", x"09", x"92", x"00", x"00", x"00", x"09", x"9C", x"00", x"00", x"00", x"09", x"A6", x"00", x"00", x"00", x"09", x"B0", x"00", x"00", x"00", x"09", x"BA", x"00", x"00", x"00", x"09", x"C4", x"00", x"00", x"00", x"09", x"CE", x"00", x"00", x"00", x"09", x"D8", x"00", x"00", x"00", x"09", x"E2", x"00", x"00", x"00", x"09", x"EC", x"00", x"00", x"00", x"09", x"F6", x"00", x"00", x"00", x"0A", x"00", x"00", x"00", x"00", x"0A", x"0A", x"00", x"00", x"00", x"0A", x"14", x"00", x"00", x"00", x"0A", x"1E", x"00", x"00", x"00", x"0A", x"28", x"00", x"00", x"00", x"0A", x"32", x"00", x"00", x"00", x"0A", x"3C", x"00", x"00", x"00", x"0A", x"46", x"00", x"00", x"00", x"0A", x"50", x"00", x"00", x"00", x"0A", x"5A", x"00", x"00", x"00", x"0A", x"64", x"00", x"00", x"00", x"0A", x"6E", x"00", x"00", x"00", x"0A", x"78", x"00", x"00", x"00", x"0A", x"82", x"00", x"00", x"00", x"0A", x"8C", x"00", x"00", x"00", x"0A", x"96", x"00", x"00", x"00", x"0A", x"A0", x"00", x"00", x"00", x"0A", x"AA", x"00", x"00", x"00", x"0A", x"B4", x"00", x"00", x"00", x"0A", x"BE", x"00", x"00", x"00", x"0A", x"C8", x"00", x"00", x"00", x"0A", x"D2", x"00", x"00", x"00", x"0A", x"DC", x"00", x"00", x"00", x"0A", x"E6", x"00", x"00", x"00", x"0A", x"F0", x"00", x"00", x"00", x"0A", x"FA", x"00", x"00", x"00", x"0B", x"04", x"00", x"00", x"00", x"0B", x"0E", x"00", x"00", x"00", x"0B", x"18", x"00", x"00", x"00", x"0B", x"22", x"00", x"00", x"00", x"0B", x"2C", x"00", x"00", x"00", x"0B", x"36", x"00", x"00", x"00", x"0B", x"40", x"00", x"00", x"00", x"0B", x"4A", x"00", x"00", x"00", x"0B", x"54", x"00", x"00", x"00", x"0B", x"5E", x"00", x"00", x"00", x"0B", x"68", x"00", x"00", x"00", x"0B", x"72", x"00", x"00", x"00", x"0B", x"7C", x"00", x"00", x"00", x"0B", x"86", x"00", x"00", x"00", x"0B", x"90", x"00", x"00", x"00", x"0B", x"9A", x"00", x"00", x"00", x"0B", x"A4", x"00", x"00", x"00", x"0B", x"AE", x"00", x"00", x"00", x"0B", x"B8", x"00", x"00", x"00", x"0B", x"C2", x"00", x"00", x"00", x"0B", x"CC", x"00", x"00", x"00", x"0B", x"D6", x"00", x"00", x"00", x"0B", x"E0", x"00", x"00", x"00", x"0B", x"EA", x"00", x"00", x"00", x"0B", x"F4", x"00", x"00", x"00", x"0B", x"FE", x"00", x"00", x"00", x"0C", x"08", x"00", x"00", x"00", x"0C", x"12", x"00", x"00", x"00", x"0C", x"1C", x"00", x"00", x"00", x"0C", x"26", x"00", x"00", x"00", x"0C", x"30", x"00", x"00", x"00", x"0C", x"3A", x"00", x"00", x"00", x"0C", x"44", x"00", x"00", x"00", x"0C", x"4E", x"00", x"00", x"00", x"0C", x"58", x"00", x"00", x"00", x"0C", x"62", x"00", x"00", x"00", x"0C", x"6C", x"00", x"00", x"00", x"0C", x"76", x"00", x"00", x"00", x"0C", x"80", x"00", x"00", x"00", x"0C", x"8A", x"00", x"00", x"00", x"0C", x"94", x"00", x"00", x"00", x"0C", x"9E", x"00", x"00", x"00", x"0C", x"A8", x"00", x"00", x"00", x"0C", x"B2", x"00", x"00", x"00", x"0C", x"BC", x"00", x"00", x"00", x"0C", x"C6", x"00", x"00", x"00", x"0C", x"D0", x"00", x"00", x"00", x"0C", x"DA", x"00", x"00", x"00", x"0C", x"E4", x"00", x"00", x"00", x"0C", x"EE", x"00", x"00", x"00", x"0C", x"F8", x"00", x"00", x"00", x"0D", x"02", x"00", x"00", x"00", x"0D", x"0C", x"00", x"00", x"00", x"0D", x"16", x"00", x"00", x"00", x"0D", x"20", x"00", x"00", x"00", x"0D", x"2A", x"00", x"00", x"00", x"0D", x"34", x"00", x"00", x"00", x"0D", x"3E", x"00", x"00", x"00", x"0D", x"48", x"00", x"00", x"00", x"0D", x"52", x"00", x"00", x"00", x"0D", x"5C", x"00", x"00", x"00", x"0D", x"66", x"00", x"00", x"00", x"0D", x"70", x"00", x"00", x"00", x"0D", x"7A", x"00", x"00", x"00", x"0D", x"84", x"00", x"00", x"00", x"0D", x"8E", x"00", x"00", x"00", x"0D", x"98", x"00", x"00", x"00", x"0D", x"A2", x"00", x"00", x"00", x"0D", x"AC", x"00", x"00", x"00", x"0D", x"B6", x"00", x"00", x"00", x"0D", x"C0", x"00", x"00", x"00", x"0D", x"CA", x"00", x"00", x"00", x"0D", x"D4", x"00", x"00", x"00", x"0D", x"DE", x"00", x"00", x"00", x"0D", x"E8", x"00", x"00", x"00", x"0D", x"F2", x"00", x"00", x"00", x"0D", x"FC", x"00", x"00", x"00", x"0E", x"06", x"00", x"00", x"00", x"0E", x"10", x"00", x"00", x"00", x"0E", x"1A", x"00", x"00", x"00", x"0E", x"24", x"00", x"00", x"00", x"0E", x"2E", x"00", x"00", x"00", x"0E", x"38", x"00", x"00", x"00", x"0E", x"42", x"00", x"00", x"00", x"0E", x"4C", x"00", x"00", x"00", x"0E", x"56", x"00", x"00", x"00", x"0E", x"60", x"00", x"00", x"00", x"0E", x"6A", x"00", x"00", x"00", x"0E", x"74", x"00", x"00", x"00", x"0E", x"7E", x"00", x"00", x"00", x"0E", x"88", x"00", x"00", x"00", x"0E", x"92", x"00", x"00", x"00", x"0E", x"9C", x"00", x"00", x"00", x"0E", x"A6", x"00", x"00", x"00", x"0E", x"B0", x"00", x"00", x"00", x"0E", x"BA", x"00", x"00", x"00", x"0E", x"C4", x"00", x"00", x"00", x"0E", x"CE", x"00", x"00", x"00", x"0E", x"D8", x"00", x"00", x"00", x"0E", x"E2", x"00", x"00", x"00", x"0E", x"EC", x"00", x"00", x"00", x"0E", x"F6", x"00", x"00", x"00", x"0F", x"00", x"00", x"00", x"00", x"0F", x"0A", x"00", x"00", x"00", x"0F", x"14", x"00", x"00", x"00", x"0F", x"1E", x"00", x"00", x"00", x"0F", x"28", x"00", x"00", x"00", x"0F", x"32", x"00", x"00", x"00", x"0F", x"3C", x"00", x"00", x"00", x"0F", x"46", x"00", x"00", x"00", x"0F", x"50", x"00", x"00", x"00", x"0F", x"5A", x"00", x"00", x"00", x"0F", x"64", x"00", x"00", x"00", x"0F", x"6E", x"00", x"00", x"00", x"0F", x"78", x"00", x"00", x"00", x"0F", x"82", x"00", x"00", x"00", x"0F", x"8C", x"00", x"00", x"00", x"0F", x"96", x"00", x"00", x"00", x"0F", x"A0", x"00", x"00", x"00", x"0F", x"AA", x"00", x"00", x"00", x"0F", x"B4", x"00", x"00", x"00", x"0F", x"BE", x"00", x"00", x"00", x"0F", x"C8", x"00", x"00", x"00", x"0F", x"D2", x"00", x"00", x"00", x"0F", x"DC", x"00", x"00", x"00", x"0F", x"E6", x"00", x"00", x"00", x"0F", x"F0", x"00", x"00", x"00", x"0F", x"FA", x"00", x"00", x"00", x"10", x"04", x"00", x"00", x"00", x"10", x"0E", x"00", x"00", x"00", x"10", x"18", x"00", x"00", x"00", x"10", x"22", x"00", x"00", x"00", x"10", x"2C", x"00", x"00", x"00", x"10", x"36", x"00", x"00", x"00", x"10", x"40", x"00", x"00", x"00", x"10", x"4A", x"00", x"00", x"00", x"10", x"54", x"00", x"00", x"00", x"10", x"5E", x"00", x"00", x"00", x"10", x"68", x"00", x"00", x"00", x"10", x"72", x"00", x"00", x"00", x"10", x"7C", x"00", x"00", x"00", x"10", x"86", x"00", x"00", x"00", x"10", x"90", x"00", x"00", x"00", x"10", x"9A", x"00", x"00", x"00", x"10", x"A4", x"00", x"00", x"00", x"10", x"AE", x"00", x"00", x"00", x"10", x"B8", x"00", x"00", x"00", x"10", x"C2", x"00", x"00", x"00", x"10", x"CC", x"00", x"00", x"00", x"10", x"D6", x"00", x"00", x"00", x"10", x"E0", x"00", x"00", x"00", x"10", x"EA", x"00", x"00", x"00", x"10", x"F4", x"00", x"00", x"00", x"10", x"FE", x"00", x"00", x"00", x"11", x"08", x"00", x"00", x"00", x"11", x"12", x"00", x"00", x"00", x"11", x"1C", x"00", x"00", x"00", x"11", x"26", x"00", x"00", x"00", x"11", x"30", x"00", x"00", x"00", x"11", x"3A", x"00", x"00", x"00", x"11", x"44", x"00", x"00", x"00", x"11", x"4E", x"00", x"00", x"00", x"11", x"58", x"00", x"00", x"00", x"11", x"62", x"00", x"00", x"00", x"11", x"6C", x"00", x"00", x"00", x"11", x"76", x"00", x"00", x"00", x"11", x"80", x"00", x"00", x"00", x"11", x"8A", x"00", x"00", x"00", x"11", x"94", x"00", x"00", x"00", x"11", x"9E", x"00", x"00", x"00", x"11", x"A8", x"00", x"00", x"00", x"11", x"B2", x"00", x"00", x"00", x"11", x"BC", x"00", x"00", x"00", x"11", x"C6", x"00", x"00", x"00", x"11", x"D0", x"00", x"00", x"00", x"11", x"DA", x"00", x"00", x"00", x"11", x"E4", x"00", x"00", x"00", x"11", x"EE", x"00", x"00", x"00", x"11", x"F8", x"00", x"00", x"00", x"12", x"02", x"00", x"00", x"00", x"12", x"0C", x"00", x"00", x"00", x"12", x"16", x"00", x"00", x"00", x"12", x"20", x"00", x"00", x"00", x"12", x"2A", x"00", x"00", x"00", x"12", x"34", x"00", x"00", x"00", x"12", x"3E", x"00", x"00", x"00", x"12", x"48", x"00", x"00", x"00", x"12", x"52", x"00", x"00", x"00", x"12", x"5C", x"00", x"00", x"00", x"12", x"66", x"00", x"00", x"00", x"12", x"70", x"00", x"00", x"00", x"12", x"7A", x"00", x"00", x"00", x"12", x"84", x"00", x"00", x"00", x"12", x"8E", x"00", x"00", x"00", x"12", x"98", x"00", x"00", x"00", x"12", x"A2", x"00", x"00", x"00", x"12", x"AC", x"00", x"00", x"00", x"12", x"B6", x"00", x"00", x"00", x"12", x"C0", x"00", x"00", x"00", x"12", x"CA", x"00", x"00", x"00", x"12", x"D4", x"00", x"00", x"00", x"12", x"DE", x"00", x"00", x"00", x"12", x"E8", x"00", x"00", x"00", x"12", x"F2", x"00", x"00", x"00", x"12", x"FC", x"00", x"00", x"00", x"13", x"06", x"00", x"00", x"00", x"13", x"10", x"00", x"00", x"00", x"13", x"1A", x"00", x"00", x"00", x"13", x"24", x"00", x"00", x"00", x"13", x"2E", x"00", x"00", x"00", x"13", x"38", x"00", x"00", x"00", x"13", x"42", x"00", x"00", x"00", x"13", x"4C", x"00", x"00", x"00", x"13", x"56", x"00", x"00", x"00", x"13", x"60", x"00", x"00", x"00", x"13", x"6A", x"00", x"00", x"00", x"13", x"74", x"00", x"00", x"00", x"13", x"7E", x"00", x"00", x"00", x"13", x"88", x"00", x"00", x"00", x"13", x"92", x"00", x"00", x"00", x"13", x"9C", x"00", x"00", x"00", x"13", x"A6", x"00", x"00", x"00", x"13", x"B0", x"00", x"00", x"00", x"13", x"BA", x"00", x"00", x"00", x"13", x"C4", x"00", x"00", x"00", x"13", x"CE", x"00", x"00", x"00", x"13", x"D8", x"00", x"00", x"00", x"13", x"E2", x"00", x"00", x"00", x"13", x"EC", x"00", x"00", x"00", x"13", x"F6", x"00", x"00", x"00", x"14", x"00", x"00", x"00", x"00", x"14", x"0A", x"00", x"00", x"00", x"14", x"14", x"00", x"00", x"00", x"14", x"1E", x"00", x"00", x"00", x"14", x"28", x"00", x"00", x"00", x"14", x"32", x"00", x"00", x"00", x"14", x"3C", x"00", x"00", x"00", x"14", x"46", x"00", x"00", x"00", x"14", x"50", x"00", x"00", x"00", x"14", x"5A", x"00", x"00", x"00", x"14", x"64", x"00", x"00", x"00", x"14", x"6E", x"00", x"00", x"00", x"14", x"78", x"00", x"00", x"00", x"14", x"82", x"00", x"00", x"00", x"14", x"8C", x"00", x"00", x"00", x"14", x"96", x"00", x"00", x"00", x"14", x"A0", x"00", x"00", x"00", x"14", x"AA", x"00", x"00", x"00", x"14", x"B4", x"00", x"00", x"00", x"14", x"BE", x"00", x"00", x"00", x"14", x"C8", x"00", x"00", x"00", x"14", x"D2", x"00", x"00", x"00", x"14", x"DC", x"00", x"00", x"00", x"14", x"E6", x"00", x"00", x"00", x"14", x"F0", x"00", x"00", x"00", x"14", x"FA", x"00", x"00", x"00", x"15", x"04", x"00", x"00", x"00", x"15", x"0E", x"00", x"00", x"00", x"15", x"18", x"00", x"00", x"00", x"15", x"22", x"00", x"00", x"00", x"15", x"2C", x"00", x"00", x"00", x"15", x"36", x"00", x"00", x"00", x"15", x"40", x"00", x"00", x"00", x"15", x"4A", x"00", x"00", x"00", x"15", x"54", x"00", x"00", x"00", x"15", x"5E", x"00", x"00", x"00", x"15", x"68", x"00", x"00", x"00", x"15", x"72", x"00", x"00", x"00", x"15", x"7C", x"00", x"00", x"00", x"15", x"86", x"00", x"00", x"00", x"15", x"90", x"00", x"00", x"00", x"15", x"9A", x"00", x"00", x"00", x"15", x"A4", x"00", x"00", x"00", x"15", x"AE", x"00", x"00", x"00", x"15", x"B8", x"00", x"00", x"00", x"15", x"C2", x"00", x"00", x"00", x"15", x"CC", x"00", x"00", x"00", x"15", x"D6", x"00", x"00", x"00", x"15", x"E0", x"00", x"00", x"00", x"15", x"EA", x"00", x"00", x"00", x"15", x"F4", x"00", x"00", x"00", x"15", x"FE", x"00", x"00", x"00", x"16", x"08", x"00", x"00", x"00", x"16", x"12", x"00", x"00", x"00", x"16", x"1C", x"00", x"00", x"00", x"16", x"26", x"00", x"00", x"00", x"16", x"30", x"00", x"00", x"00", x"16", x"3A", x"00", x"00", x"00", x"16", x"44", x"00", x"00", x"00", x"16", x"4E", x"00", x"00", x"00", x"16", x"58", x"00", x"00", x"00", x"16", x"62", x"00", x"00", x"00", x"16", x"6C", x"00", x"00", x"00", x"16", x"76", x"00", x"00", x"00", x"16", x"80", x"00", x"00", x"00", x"16", x"8A", x"00", x"00", x"00", x"16", x"94", x"00", x"00", x"00", x"16", x"9E", x"00", x"00", x"00", x"16", x"A8", x"00", x"00", x"00", x"16", x"B2", x"00", x"00", x"00", x"16", x"BC", x"00", x"00", x"00", x"16", x"C6", x"00", x"00", x"00", x"16", x"D0", x"00", x"00", x"00", x"16", x"DA", x"00", x"00", x"00", x"16", x"E4", x"00", x"00", x"00", x"16", x"EE", x"00", x"00", x"00", x"16", x"F8", x"00", x"00", x"00", x"17", x"02", x"00", x"00", x"00", x"17", x"0C", x"00", x"00", x"00", x"17", x"16", x"00", x"00", x"00", x"17", x"20", x"00", x"00", x"00", x"17", x"2A", x"00", x"00", x"00", x"17", x"34", x"00", x"00", x"00", x"17", x"3E", x"00", x"00", x"00", x"17", x"48", x"00", x"00", x"00", x"17", x"52", x"00", x"00", x"00", x"17", x"5C", x"00", x"00", x"00", x"17", x"66", x"00", x"00", x"00", x"17", x"70", x"00", x"00", x"00", x"17", x"7A", x"00", x"00", x"00", x"17", x"84", x"00", x"00", x"00", x"17", x"8E", x"00", x"00", x"00", x"17", x"98", x"00", x"00", x"00", x"17", x"A2", x"00", x"00", x"00", x"17", x"AC", x"00", x"00", x"00", x"17", x"B6", x"00", x"00", x"00", x"17", x"C0", x"00", x"00", x"00", x"17", x"CA", x"00", x"00", x"00", x"17", x"D4", x"00", x"00", x"00", x"17", x"DE", x"00", x"00", x"00", x"17", x"E8", x"00", x"00", x"00", x"17", x"F2", x"00", x"00", x"00", x"17", x"FC", x"00", x"00", x"00", x"18", x"06", x"00", x"00", x"00", x"18", x"10", x"00", x"00", x"00", x"18", x"1A", x"00", x"00", x"00", x"18", x"24", x"00", x"00", x"00", x"18", x"2E", x"00", x"00", x"00", x"18", x"38", x"00", x"00", x"00", x"18", x"42", x"00", x"00", x"00", x"18", x"4C", x"00", x"00", x"00", x"18", x"56", x"00", x"00", x"00", x"18", x"60", x"00", x"00", x"00", x"18", x"6A", x"00", x"00", x"00", x"18", x"74", x"00", x"00", x"00", x"18", x"7E", x"00", x"00", x"00", x"18", x"88", x"00", x"00", x"00", x"18", x"92", x"00", x"00", x"00", x"18", x"9C", x"00", x"00", x"00", x"18", x"A6", x"00", x"00", x"00", x"18", x"B0", x"00", x"00", x"00", x"18", x"BA", x"00", x"00", x"00", x"18", x"C4", x"00", x"00", x"00", x"18", x"CE", x"00", x"00", x"00", x"18", x"D8", x"00", x"00", x"00", x"18", x"E2", x"00", x"00", x"00", x"18", x"EC", x"00", x"00", x"00", x"18", x"F6", x"00", x"00", x"00", x"19", x"00", x"00", x"00", x"00", x"19", x"0A", x"00", x"00", x"00", x"19", x"14", x"00", x"00", x"00", x"19", x"1E", x"00", x"00", x"00", x"19", x"28", x"00", x"00", x"00", x"19", x"32", x"00", x"00", x"00", x"19", x"3C", x"00", x"00", x"00", x"19", x"46", x"00", x"00", x"00", x"19", x"50", x"00", x"00", x"00", x"19", x"5A", x"00", x"00", x"00", x"19", x"64", x"00", x"00", x"00", x"19", x"6E", x"00", x"00", x"00", x"19", x"78", x"00", x"00", x"00", x"19", x"82", x"00", x"00", x"00", x"19", x"8C", x"00", x"00", x"00", x"19", x"96", x"00", x"00", x"00", x"19", x"A0", x"00", x"00", x"00", x"19", x"AA", x"00", x"00", x"00", x"19", x"B4", x"00", x"00", x"00", x"19", x"BE", x"00", x"00", x"00", x"19", x"C8", x"00", x"00", x"00", x"19", x"D2", x"00", x"00", x"00", x"19", x"DC", x"00", x"00", x"00", x"19", x"E6", x"00", x"00", x"00", x"19", x"F0", x"00", x"00", x"00", x"19", x"FA", x"00", x"00", x"00", x"1A", x"04", x"00", x"00", x"00", x"1A", x"0E", x"00", x"00", x"00", x"1A", x"18", x"00", x"00", x"00", x"1A", x"22", x"00", x"00", x"00", x"1A", x"2C", x"00", x"00", x"00", x"1A", x"36", x"00", x"00", x"00", x"1A", x"40", x"00", x"00", x"00", x"1A", x"4A", x"00", x"00", x"00", x"1A", x"54", x"00", x"00", x"00", x"1A", x"5E", x"00", x"00", x"00", x"1A", x"68", x"00", x"00", x"00", x"1A", x"72", x"00", x"00", x"00", x"1A", x"7C", x"00", x"00", x"00", x"1A", x"86", x"00", x"00", x"00", x"1A", x"90", x"00", x"00", x"00", x"1A", x"9A", x"00", x"00", x"00", x"1A", x"A4", x"00", x"00", x"00", x"1A", x"AE", x"00", x"00", x"00", x"1A", x"B8", x"00", x"00", x"00", x"1A", x"C2", x"00", x"00", x"00", x"1A", x"CC", x"00", x"00", x"00", x"1A", x"D6", x"00", x"00", x"00", x"1A", x"E0", x"00", x"00", x"00", x"1A", x"EA", x"00", x"00", x"00", x"1A", x"F4", x"00", x"00", x"00", x"1A", x"FE", x"00", x"00", x"00", x"1B", x"08", x"00", x"00", x"00", x"1B", x"12", x"00", x"00", x"00", x"1B", x"1C", x"00", x"00", x"00", x"1B", x"26", x"00", x"00", x"00", x"1B", x"30", x"00", x"00", x"00", x"1B", x"3A", x"00", x"00", x"00", x"1B", x"44", x"00", x"00", x"00", x"1B", x"4E", x"00", x"00", x"00", x"1B", x"58", x"00", x"00", x"00", x"1B", x"62", x"00", x"00", x"00", x"1B", x"6C", x"00", x"00", x"00", x"1B", x"76", x"00", x"00", x"00", x"1B", x"80", x"00", x"00", x"00", x"1B", x"8A", x"00", x"00", x"00", x"1B", x"94", x"00", x"00", x"00", x"1B", x"9E", x"00", x"00", x"00", x"1B", x"A8", x"00", x"00", x"00", x"1B", x"B2", x"00", x"00", x"00", x"1B", x"BC", x"00", x"00", x"00", x"1B", x"C6", x"00", x"00", x"00", x"1B", x"D0", x"00", x"00", x"00", x"1B", x"DA", x"00", x"00", x"00", x"1B", x"E4", x"00", x"00", x"00", x"1B", x"EE", x"00", x"00", x"00", x"1B", x"F8", x"00", x"00", x"00", x"1C", x"02", x"00", x"00", x"00", x"1C", x"0C", x"00", x"00", x"00", x"1C", x"16", x"00", x"00", x"00", x"1C", x"20", x"00", x"00", x"00", x"1C", x"2A", x"00", x"00", x"00", x"1C", x"34", x"00", x"00", x"00", x"1C", x"3E", x"00", x"00", x"00", x"1C", x"48", x"00", x"00", x"00", x"1C", x"52", x"00", x"00", x"00", x"1C", x"5C", x"00", x"00", x"00", x"1C", x"66", x"00", x"00", x"00", x"1C", x"70", x"00", x"00", x"00", x"1C", x"7A", x"00", x"00", x"00", x"1C", x"84", x"00", x"00", x"00", x"1C", x"8E", x"00", x"00", x"00", x"1C", x"98", x"00", x"00", x"00", x"1C", x"A2", x"00", x"00", x"00", x"1C", x"AC", x"00", x"00", x"00", x"1C", x"B6", x"00", x"00", x"00", x"1C", x"C0", x"00", x"00", x"00", x"1C", x"CA", x"00", x"00", x"00", x"1C", x"D4", x"00", x"00", x"00", x"1C", x"DE", x"00", x"00", x"00", x"1C", x"E8", x"00", x"00", x"00", x"1C", x"F2", x"00", x"00", x"00", x"1C", x"FC", x"00", x"00", x"00", x"1D", x"06", x"00", x"00", x"00", x"1D", x"10", x"00", x"00", x"00", x"1D", x"1A", x"00", x"00", x"00", x"1D", x"24", x"00", x"00", x"00", x"1D", x"2E", x"00", x"00", x"00", x"1D", x"38", x"00", x"00", x"00", x"1D", x"42", x"00", x"00", x"00", x"1D", x"4C", x"00", x"00", x"00", x"1D", x"56", x"00", x"00", x"00", x"1D", x"60", x"00", x"00", x"00", x"1D", x"6A", x"00", x"00", x"00", x"1D", x"74", x"00", x"00", x"00", x"1D", x"7E", x"00", x"00", x"00", x"1D", x"88", x"00", x"00", x"00", x"1D", x"92", x"00", x"00", x"00", x"1D", x"9C", x"00", x"00", x"00", x"1D", x"A6", x"00", x"00", x"00", x"1D", x"B0", x"00", x"00", x"00", x"1D", x"BA", x"00", x"00", x"00", x"1D", x"C4", x"00", x"00", x"00", x"1D", x"CE", x"00", x"00", x"00", x"1D", x"D8", x"00", x"00", x"00", x"1D", x"E2", x"00", x"00", x"00", x"1D", x"EC", x"00", x"00", x"00", x"1D", x"F6", x"00", x"00", x"00", x"1E", x"00", x"00", x"00", x"00", x"1E", x"0A", x"00", x"00", x"00", x"1E", x"14", x"00", x"00", x"00", x"1E", x"1E", x"00", x"00", x"00", x"1E", x"28", x"00", x"00", x"00", x"1E", x"32", x"00", x"00", x"00", x"1E", x"3C", x"00", x"00", x"00", x"1E", x"46", x"00", x"00", x"00", x"1E", x"50", x"00", x"00", x"00", x"1E", x"5A", x"00", x"00", x"00", x"1E", x"64", x"00", x"00", x"00", x"1E", x"6E", x"00", x"00", x"00", x"1E", x"78", x"00", x"00", x"00", x"1E", x"82", x"00", x"00", x"00", x"1E", x"8C", x"00", x"00", x"00", x"1E", x"96", x"00", x"00", x"00", x"1E", x"A0", x"00", x"00", x"00", x"1E", x"AA", x"00", x"00", x"00", x"1E", x"B4", x"00", x"00", x"00", x"1E", x"BE", x"00", x"00", x"00", x"1E", x"C8", x"00", x"00", x"00", x"1E", x"D2", x"00", x"00", x"00", x"1E", x"DC", x"00", x"00", x"00", x"1E", x"E6", x"00", x"00", x"00", x"1E", x"F0", x"00", x"00", x"00", x"1E", x"FA", x"00", x"00", x"00", x"1F", x"04", x"00", x"00", x"00", x"1F", x"0E", x"00", x"00", x"00", x"1F", x"18", x"00", x"00", x"00", x"1F", x"22", x"00", x"00", x"00", x"1F", x"2C", x"00", x"00", x"00", x"1F", x"36", x"00", x"00", x"00", x"1F", x"40", x"00", x"00", x"00", x"1F", x"4A", x"00", x"00", x"00", x"1F", x"54", x"00", x"00", x"00", x"1F", x"5E", x"00", x"00", x"00", x"1F", x"68", x"00", x"00", x"00", x"1F", x"72", x"00", x"00", x"00", x"1F", x"7C", x"00", x"00", x"00", x"1F", x"86", x"00", x"00", x"00", x"1F", x"90", x"00", x"00", x"00", x"1F", x"9A", x"00", x"00", x"00", x"1F", x"A4", x"00", x"00", x"00", x"1F", x"AE", x"00", x"00", x"00", x"1F", x"B8", x"00", x"00", x"00", x"1F", x"C2", x"00", x"00", x"00", x"1F", x"CC", x"00", x"00", x"00", x"1F", x"D6", x"00", x"00", x"00", x"1F", x"E0", x"00", x"00", x"00", x"1F", x"EA", x"00", x"00", x"00", x"1F", x"F4", x"00", x"00", x"00", x"1F", x"FE", x"00", x"00", x"00", x"20", x"08", x"00", x"00", x"00", x"20", x"12", x"00", x"00", x"00", x"20", x"1C", x"00", x"00", x"00", x"20", x"26", x"00", x"00", x"00", x"20", x"30", x"00", x"00", x"00", x"20", x"3A", x"00", x"00", x"00", x"20", x"44", x"00", x"00", x"00", x"20", x"4E", x"00", x"00", x"00", x"20", x"58", x"00", x"00", x"00", x"20", x"62", x"00", x"00", x"00", x"20", x"6C", x"00", x"00", x"00", x"20", x"76", x"00", x"00", x"00", x"20", x"80", x"00", x"00", x"00", x"20", x"8A", x"00", x"00", x"00", x"20", x"94", x"00", x"00", x"00", x"20", x"9E", x"00", x"00", x"00", x"20", x"A8", x"00", x"00", x"00", x"20", x"B2", x"00", x"00", x"00", x"20", x"BC", x"00", x"00", x"00", x"20", x"C6", x"00", x"00", x"00", x"20", x"D0", x"00", x"00", x"00", x"20", x"DA", x"00", x"00", x"00", x"20", x"E4", x"00", x"00", x"00", x"20", x"EE", x"00", x"00", x"00", x"20", x"F8", x"00", x"00", x"00", x"21", x"02", x"00", x"00", x"00", x"21", x"0C", x"00", x"00", x"00", x"21", x"16", x"00", x"00", x"00", x"21", x"20", x"00", x"00", x"00", x"21", x"2A", x"00", x"00", x"00", x"21", x"34", x"00", x"00", x"00", x"21", x"3E", x"00", x"00", x"00", x"21", x"48", x"00", x"00", x"00", x"21", x"52", x"00", x"00", x"00", x"21", x"5C", x"00", x"00", x"00", x"21", x"66", x"00", x"00", x"00", x"21", x"70", x"00", x"00", x"00", x"21", x"7A", x"00", x"00", x"00", x"21", x"84", x"00", x"00", x"00", x"21", x"8E", x"00", x"00", x"00", x"21", x"98", x"00", x"00", x"00", x"21", x"A2", x"00", x"00", x"00", x"21", x"AC", x"00", x"00", x"00", x"21", x"B6", x"00", x"00", x"00", x"21", x"C0", x"00", x"00", x"00", x"21", x"CA", x"00", x"00", x"00", x"21", x"D4", x"00", x"00", x"00", x"21", x"DE", x"00", x"00", x"00", x"21", x"E8", x"00", x"00", x"00", x"21", x"F2", x"00", x"00", x"00", x"21", x"FC", x"00", x"00", x"00", x"22", x"06", x"00", x"00", x"00", x"22", x"10", x"00", x"00", x"00", x"22", x"1A", x"00", x"00", x"00", x"22", x"24", x"00", x"00", x"00", x"22", x"2E", x"00", x"00", x"00", x"22", x"38", x"00", x"00", x"00", x"22", x"42", x"00", x"00", x"00", x"22", x"4C", x"00", x"00", x"00", x"22", x"56", x"00", x"00", x"00", x"22", x"60", x"00", x"00", x"00", x"22", x"6A", x"00", x"00", x"00", x"22", x"74", x"00", x"00", x"00", x"22", x"7E", x"00", x"00", x"00", x"22", x"88", x"00", x"00", x"00", x"22", x"92", x"00", x"00", x"00", x"22", x"9C", x"00", x"00", x"00", x"22", x"A6", x"00", x"00", x"00", x"22", x"B0", x"00", x"00", x"00", x"22", x"BA", x"00", x"00", x"00", x"22", x"C4", x"00", x"00", x"00", x"22", x"CE", x"00", x"00", x"00", x"22", x"D8", x"00", x"00", x"00", x"22", x"E2", x"00", x"00", x"00", x"22", x"EC", x"00", x"00", x"00", x"22", x"F6", x"00", x"00", x"00", x"23", x"00", x"00", x"00", x"00", x"23", x"0A", x"00", x"00", x"00", x"23", x"14", x"00", x"00", x"00", x"23", x"1E", x"00", x"00", x"00", x"23", x"28", x"00", x"00", x"00", x"23", x"32", x"00", x"00", x"00", x"23", x"3C", x"00", x"00", x"00", x"23", x"46", x"00", x"00", x"00", x"23", x"50", x"00", x"00", x"00", x"23", x"5A", x"00", x"00", x"00", x"23", x"64", x"00", x"00", x"00", x"23", x"6E", x"00", x"00", x"00", x"23", x"78", x"00", x"00", x"00", x"23", x"82", x"00", x"00", x"00", x"23", x"8C", x"00", x"00", x"00", x"23", x"96", x"00", x"00", x"00", x"23", x"A0", x"00", x"00", x"00", x"23", x"AA", x"00", x"00", x"00", x"23", x"B4", x"00", x"00", x"00", x"23", x"BE", x"00", x"00", x"00", x"23", x"C8", x"00", x"00", x"00", x"23", x"D2", x"00", x"00", x"00", x"23", x"DC", x"00", x"00", x"00", x"23", x"E6", x"00", x"00", x"00", x"23", x"F0", x"00", x"00", x"00", x"23", x"FA", x"00", x"00", x"00", x"24", x"04", x"00", x"00", x"00", x"24", x"0E", x"00", x"00", x"00", x"24", x"18", x"00", x"00", x"00", x"24", x"22", x"00", x"00", x"00", x"24", x"2C", x"00", x"00", x"00", x"24", x"36", x"00", x"00", x"00", x"24", x"40", x"00", x"00", x"00", x"24", x"4A", x"00", x"00", x"00", x"24", x"54", x"00", x"00", x"00", x"24", x"5E", x"00", x"00", x"00", x"24", x"68", x"00", x"00", x"00", x"24", x"72", x"00", x"00", x"00", x"24", x"7C", x"00", x"00", x"00", x"24", x"86", x"00", x"00", x"00", x"24", x"90", x"00", x"00", x"00", x"24", x"9A", x"00", x"00", x"00", x"24", x"A4", x"00", x"00", x"00", x"24", x"AE", x"00", x"00", x"00", x"24", x"B8", x"00", x"00", x"00", x"24", x"C2", x"00", x"00", x"00", x"24", x"CC", x"00", x"00", x"00", x"24", x"D6", x"00", x"00", x"00", x"24", x"E0", x"00", x"00", x"00", x"24", x"EA", x"00", x"00", x"00", x"24", x"F4", x"00", x"00", x"00", x"24", x"FE", x"00", x"00", x"00", x"25", x"08", x"00", x"00", x"00", x"25", x"12", x"00", x"00", x"00", x"25", x"1C", x"00", x"00", x"00", x"25", x"26", x"00", x"00", x"00", x"25", x"30", x"00", x"00", x"00", x"25", x"3A", x"00", x"00", x"00", x"25", x"44", x"00", x"00", x"00", x"25", x"4E", x"00", x"00", x"00", x"25", x"58", x"00", x"00", x"00", x"25", x"62", x"00", x"00", x"00", x"25", x"6C", x"00", x"00", x"00", x"25", x"76", x"00", x"00", x"00", x"25", x"80", x"00", x"00", x"00", x"25", x"8A", x"00", x"00", x"00", x"25", x"94", x"00", x"00", x"00", x"25", x"9E", x"00", x"00", x"00", x"25", x"A8", x"00", x"00", x"00", x"25", x"B2", x"00", x"00", x"00", x"25", x"BC", x"00", x"00", x"00", x"25", x"C6", x"00", x"00", x"00", x"25", x"D0", x"00", x"00", x"00", x"25", x"DA", x"00", x"00", x"00", x"25", x"E4", x"00", x"00", x"00", x"25", x"EE", x"00", x"00", x"00", x"25", x"F8", x"00", x"00", x"00", x"26", x"02", x"00", x"00", x"00", x"26", x"0C", x"00", x"00", x"00", x"26", x"16", x"00", x"00", x"00", x"26", x"20", x"00", x"00", x"00", x"26", x"2A", x"00", x"00", x"00", x"26", x"34", x"00", x"00", x"00", x"26", x"3E", x"00", x"00", x"00", x"26", x"48", x"00", x"00", x"00", x"26", x"52", x"00", x"00", x"00", x"26", x"5C", x"00", x"00", x"00", x"26", x"66", x"00", x"00", x"00", x"26", x"70", x"00", x"00", x"00", x"26", x"7A", x"00", x"00", x"00", x"26", x"84", x"00", x"00", x"00", x"26", x"8E", x"00", x"00", x"00", x"26", x"98", x"00", x"00", x"00", x"26", x"A2", x"00", x"00", x"00", x"26", x"AC", x"00", x"00", x"00", x"26", x"B6", x"00", x"00", x"00", x"26", x"C0", x"00", x"00", x"00", x"26", x"CA", x"00", x"00", x"00", x"26", x"D4", x"00", x"00", x"00", x"26", x"DE", x"00", x"00", x"00", x"26", x"E8", x"00", x"00", x"00", x"26", x"F2", x"00", x"00", x"00", x"26", x"FC", x"00", x"00", x"00", x"27", x"06", x"00", x"00", x"00", x"27", x"10", x"00", x"00", x"00", x"27", x"1A", x"00", x"00", x"00", x"27", x"24", x"00", x"00", x"00", x"27", x"2E", x"00", x"00", x"00", x"27", x"38", x"00", x"00", x"00", x"27", x"42", x"00", x"00", x"00", x"27", x"4C", x"00", x"00", x"00", x"27", x"56", x"00", x"00", x"00", x"27", x"60", x"00", x"00", x"00", x"27", x"6A", x"00", x"00", x"00", x"27", x"74", x"00", x"00", x"00", x"27", x"7E", x"00", x"00", x"00", x"27", x"88", x"00", x"00", x"00", x"27", x"92", x"00", x"00", x"00", x"27", x"9C", x"00", x"00", x"00", x"27", x"A6", x"00", x"00", x"00", x"27", x"B0", x"00", x"00", x"00", x"27", x"BA", x"00", x"00", x"00", x"27", x"C4", x"00", x"00", x"00", x"27", x"CE", x"00", x"00", x"00", x"27", x"D8", x"00", x"00", x"00", x"27", x"E2", x"00", x"00", x"00", x"27", x"EC", x"00", x"00", x"00", x"27", x"F6", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"0A", x"00", x"00", x"00", x"00", x"14", x"00", x"00", x"00", x"00", x"1E", x"00", x"00", x"00", x"00", x"28", x"00", x"00", x"00", x"00", x"32", x"00", x"00", x"00", x"00", x"3C", x"00", x"00", x"00", x"00", x"46", x"00", x"00", x"00", x"00", x"50", x"00", x"00", x"00", x"00", x"5A", x"00", x"00", x"00", x"00", x"64", x"00", x"00", x"00", x"00", x"6E", x"00", x"00", x"00", x"00", x"78", x"00", x"00", x"00", x"00", x"82", x"00", x"00", x"00", x"00", x"8C", x"00", x"00", x"00", x"00", x"96", x"00", x"00", x"00", x"00", x"A0", x"00", x"00", x"00", x"00", x"AA", x"00", x"00", x"00", x"00", x"B4", x"00", x"00", x"00", x"00", x"BE", x"00", x"00", x"00", x"00", x"C8", x"00", x"00", x"00", x"00", x"D2", x"00", x"00", x"00", x"00", x"DC", x"00", x"00", x"00", x"00", x"E6", x"00", x"00", x"00", x"00", x"F0", x"00", x"00", x"00", x"00", x"FA", x"00", x"00", x"00", x"01", x"04", x"00", x"00", x"00", x"01", x"0E", x"00", x"00", x"00", x"01", x"18", x"00", x"00", x"00", x"01", x"22", x"00", x"00", x"00", x"01", x"2C", x"00", x"00", x"00", x"01", x"36", x"00", x"00", x"00", x"01", x"40", x"00", x"00", x"00", x"01", x"4A", x"00", x"00", x"00", x"01", x"54", x"00", x"00", x"00", x"01", x"5E", x"00", x"00", x"00", x"01", x"68", x"00", x"00", x"00", x"01", x"72", x"00", x"00", x"00", x"01", x"7C", x"00", x"00", x"00", x"01", x"86", x"00", x"00", x"00", x"01", x"90", x"00", x"00", x"00", x"01", x"9A", x"00", x"00", x"00", x"01", x"A4", x"00", x"00", x"00", x"01", x"AE", x"00", x"00", x"00", x"01", x"B8", x"00", x"00", x"00", x"01", x"C2", x"00", x"00", x"00", x"01", x"CC", x"00", x"00", x"00", x"01", x"D6", x"00", x"00", x"00", x"01", x"E0", x"00", x"00", x"00", x"01", x"EA", x"00", x"00", x"00", x"01", x"F4", x"00", x"00", x"00", x"01", x"FE", x"00", x"00", x"00", x"02", x"08", x"00", x"00", x"00", x"02", x"12", x"00", x"00", x"00", x"02", x"1C", x"00", x"00", x"00", x"02", x"26", x"00", x"00", x"00", x"02", x"30", x"00", x"00", x"00", x"02", x"3A", x"00", x"00", x"00", x"02", x"44", x"00", x"00", x"00", x"02", x"4E", x"00", x"00", x"00", x"02", x"58", x"00", x"00", x"00", x"02", x"62", x"00", x"00", x"00", x"02", x"6C", x"00", x"00", x"00", x"02", x"76", x"00", x"00", x"00", x"02", x"80", x"00", x"00", x"00", x"02", x"8A", x"00", x"00", x"00", x"02", x"94", x"00", x"00", x"00", x"02", x"9E", x"00", x"00", x"00", x"02", x"A8", x"00", x"00", x"00", x"02", x"B2", x"00", x"00", x"00", x"02", x"BC", x"00", x"00", x"00", x"02", x"C6", x"00", x"00", x"00", x"02", x"D0", x"00", x"00", x"00", x"02", x"DA", x"00", x"00", x"00", x"02", x"E4", x"00", x"00", x"00", x"02", x"EE", x"00", x"00", x"00", x"02", x"F8", x"00", x"00", x"00", x"03", x"02", x"00", x"00", x"00", x"03", x"0C", x"00", x"00", x"00", x"03", x"16", x"00", x"00", x"00", x"03", x"20", x"00", x"00", x"00", x"03", x"2A", x"00", x"00", x"00", x"03", x"34", x"00", x"00", x"00", x"03", x"3E", x"00", x"00", x"00", x"03", x"48", x"00", x"00", x"00", x"03", x"52", x"00", x"00", x"00", x"03", x"5C", x"00", x"00", x"00", x"03", x"66", x"00", x"00", x"00", x"03", x"70", x"00", x"00", x"00", x"03", x"7A", x"00", x"00", x"00", x"03", x"84", x"00", x"00", x"00", x"03", x"8E", x"00", x"00", x"00", x"03", x"98", x"00", x"00", x"00", x"03", x"A2", x"00", x"00", x"00", x"03", x"AC", x"00", x"00", x"00", x"03", x"B6", x"00", x"00", x"00", x"03", x"C0", x"00", x"00", x"00", x"03", x"CA", x"00", x"00", x"00", x"03", x"D4", x"00", x"00", x"00", x"03", x"DE", x"00", x"00", x"00", x"03", x"E8", x"00", x"00", x"00", x"03", x"F2", x"00", x"00", x"00", x"03", x"FC", x"00", x"00", x"00", x"04", x"06", x"00", x"00", x"00", x"04", x"10", x"00", x"00", x"00", x"04", x"1A", x"00", x"00", x"00", x"04", x"24", x"00", x"00", x"00", x"04", x"2E", x"00", x"00", x"00", x"04", x"38", x"00", x"00", x"00", x"04", x"42", x"00", x"00", x"00", x"04", x"4C", x"00", x"00", x"00", x"04", x"56", x"00", x"00", x"00", x"04", x"60", x"00", x"00", x"00", x"04", x"6A", x"00", x"00", x"00", x"04", x"74", x"00", x"00", x"00", x"04", x"7E", x"00", x"00", x"00", x"04", x"88", x"00", x"00", x"00", x"04", x"92", x"00", x"00", x"00", x"04", x"9C", x"00", x"00", x"00", x"04", x"A6", x"00", x"00", x"00", x"04", x"B0", x"00", x"00", x"00", x"04", x"BA", x"00", x"00", x"00", x"04", x"C4", x"00", x"00", x"00", x"04", x"CE", x"00", x"00", x"00", x"04", x"D8", x"00", x"00", x"00", x"04", x"E2", x"00", x"00", x"00", x"04", x"EC", x"00", x"00", x"00", x"04", x"F6", x"00", x"00", x"00", x"05", x"00", x"00", x"00", x"00", x"05", x"0A", x"00", x"00", x"00", x"05", x"14", x"00", x"00", x"00", x"05", x"1E", x"00", x"00", x"00", x"05", x"28", x"00", x"00", x"00", x"05", x"32", x"00", x"00", x"00", x"05", x"3C", x"00", x"00", x"00", x"05", x"46", x"00", x"00", x"00", x"05", x"50", x"00", x"00", x"00", x"05", x"5A", x"00", x"00", x"00", x"05", x"64", x"00", x"00", x"00", x"05", x"6E", x"00", x"00", x"00", x"05", x"78", x"00", x"00", x"00", x"05", x"82", x"00", x"00", x"00", x"05", x"8C", x"00", x"00", x"00", x"05", x"96", x"00", x"00", x"00", x"05", x"A0", x"00", x"00", x"00", x"05", x"AA", x"00", x"00", x"00", x"05", x"B4", x"00", x"00", x"00", x"05", x"BE", x"00", x"00", x"00", x"05", x"C8", x"00", x"00", x"00", x"05", x"D2", x"00", x"00", x"00", x"05", x"DC", x"00", x"00", x"00", x"05", x"E6", x"00", x"00", x"00", x"05", x"F0", x"00", x"00", x"00", x"05", x"FA", x"00", x"00", x"00", x"06", x"04", x"00", x"00", x"00", x"06", x"0E", x"00", x"00", x"00", x"06", x"18", x"00", x"00", x"00", x"06", x"22", x"00", x"00", x"00", x"06", x"2C", x"00", x"00", x"00", x"06", x"36", x"00", x"00", x"00", x"06", x"40", x"00", x"00", x"00", x"06", x"4A", x"00", x"00", x"00", x"06", x"54", x"00", x"00", x"00", x"06", x"5E", x"00", x"00", x"00", x"06", x"68", x"00", x"00", x"00", x"06", x"72", x"00", x"00", x"00", x"06", x"7C", x"00", x"00", x"00", x"06", x"86", x"00", x"00", x"00", x"06", x"90", x"00", x"00", x"00", x"06", x"9A", x"00", x"00", x"00", x"06", x"A4", x"00", x"00", x"00", x"06", x"AE", x"00", x"00", x"00", x"06", x"B8", x"00", x"00", x"00", x"06", x"C2", x"00", x"00", x"00", x"06", x"CC", x"00", x"00", x"00", x"06", x"D6", x"00", x"00", x"00", x"06", x"E0", x"00", x"00", x"00", x"06", x"EA", x"00", x"00", x"00", x"06", x"F4", x"00", x"00", x"00", x"06", x"FE", x"00", x"00", x"00", x"07", x"08", x"00", x"00", x"00", x"07", x"12", x"00", x"00", x"00", x"07", x"1C", x"00", x"00", x"00", x"07", x"26", x"00", x"00", x"00", x"07", x"30", x"00", x"00", x"00", x"07", x"3A", x"00", x"00", x"00", x"07", x"44", x"00", x"00", x"00", x"07", x"4E", x"00", x"00", x"00", x"07", x"58", x"00", x"00", x"00", x"07", x"62", x"00", x"00", x"00", x"07", x"6C", x"00", x"00", x"00", x"07", x"76", x"00", x"00", x"00", x"07", x"80", x"00", x"00", x"00", x"07", x"8A", x"00", x"00", x"00", x"07", x"94", x"00", x"00", x"00", x"07", x"9E", x"00", x"00", x"00", x"07", x"A8", x"00", x"00", x"00", x"07", x"B2", x"00", x"00", x"00", x"07", x"BC", x"00", x"00", x"00", x"07", x"C6", x"00", x"00", x"00", x"07", x"D0", x"00", x"00", x"00", x"07", x"DA", x"00", x"00", x"00", x"07", x"E4", x"00", x"00", x"00", x"07", x"EE", x"00", x"00", x"00", x"07", x"F8", x"00", x"00", x"00", x"08", x"02", x"00", x"00", x"00", x"08", x"0C", x"00", x"00", x"00", x"08", x"16", x"00", x"00", x"00", x"08", x"20", x"00", x"00", x"00", x"08", x"2A", x"00", x"00", x"00", x"08", x"34", x"00", x"00", x"00", x"08", x"3E", x"00", x"00", x"00", x"08", x"48", x"00", x"00", x"00", x"08", x"52", x"00", x"00", x"00", x"08", x"5C", x"00", x"00", x"00", x"08", x"66", x"00", x"00", x"00", x"08", x"70", x"00", x"00", x"00", x"08", x"7A", x"00", x"00", x"00", x"08", x"84", x"00", x"00", x"00", x"08", x"8E", x"00", x"00", x"00", x"08", x"98", x"00", x"00", x"00", x"08", x"A2", x"00", x"00", x"00", x"08", x"AC", x"00", x"00", x"00", x"08", x"B6", x"00", x"00", x"00", x"08", x"C0", x"00", x"00", x"00", x"08", x"CA", x"00", x"00", x"00", x"08", x"D4", x"00", x"00", x"00", x"08", x"DE", x"00", x"00", x"00", x"08", x"E8", x"00", x"00", x"00", x"08", x"F2", x"00", x"00", x"00", x"08", x"FC", x"00", x"00", x"00", x"09", x"06", x"00", x"00", x"00", x"09", x"10", x"00", x"00", x"00", x"09", x"1A", x"00", x"00", x"00", x"09", x"24", x"00", x"00", x"00", x"09", x"2E", x"00", x"00", x"00", x"09", x"38", x"00", x"00", x"00", x"09", x"42", x"00", x"00", x"00", x"09", x"4C", x"00", x"00", x"00", x"09", x"56", x"00", x"00", x"00", x"09", x"60", x"00", x"00", x"00", x"09", x"6A", x"00", x"00", x"00", x"09", x"74", x"00", x"00", x"00", x"09", x"7E", x"00", x"00", x"00", x"09", x"88", x"00", x"00", x"00", x"09", x"92", x"00", x"00", x"00", x"09", x"9C", x"00", x"00", x"00", x"09", x"A6", x"00", x"00", x"00", x"09", x"B0", x"00", x"00", x"00", x"09", x"BA", x"00", x"00", x"00", x"09", x"C4", x"00", x"00", x"00", x"09", x"CE", x"00", x"00", x"00", x"09", x"D8", x"00", x"00", x"00", x"09", x"E2", x"00", x"00", x"00", x"09", x"EC", x"00", x"00", x"00", x"09", x"F6", x"00", x"00", x"00", x"0A", x"00", x"00", x"00", x"00", x"0A", x"0A", x"00", x"00", x"00", x"0A", x"14", x"00", x"00", x"00", x"0A", x"1E", x"00", x"00", x"00", x"0A", x"28", x"00", x"00", x"00", x"0A", x"32", x"00", x"00", x"00", x"0A", x"3C", x"00", x"00", x"00", x"0A", x"46", x"00", x"00", x"00", x"0A", x"50", x"00", x"00", x"00", x"0A", x"5A", x"00", x"00", x"00", x"0A", x"64", x"00", x"00", x"00", x"0A", x"6E", x"00", x"00", x"00", x"0A", x"78", x"00", x"00", x"00", x"0A", x"82", x"00", x"00", x"00", x"0A", x"8C", x"00", x"00", x"00", x"0A", x"96", x"00", x"00", x"00", x"0A", x"A0", x"00", x"00", x"00", x"0A", x"AA", x"00", x"00", x"00", x"0A", x"B4", x"00", x"00", x"00", x"0A", x"BE", x"00", x"00", x"00", x"0A", x"C8", x"00", x"00", x"00", x"0A", x"D2", x"00", x"00", x"00", x"0A", x"DC", x"00", x"00", x"00", x"0A", x"E6", x"00", x"00", x"00", x"0A", x"F0", x"00", x"00", x"00", x"0A", x"FA", x"00", x"00", x"00", x"0B", x"04", x"00", x"00", x"00", x"0B", x"0E", x"00", x"00", x"00", x"0B", x"18", x"00", x"00", x"00", x"0B", x"22", x"00", x"00", x"00", x"0B", x"2C", x"00", x"00", x"00", x"0B", x"36", x"00", x"00", x"00", x"0B", x"40", x"00", x"00", x"00", x"0B", x"4A", x"00", x"00", x"00", x"0B", x"54", x"00", x"00", x"00", x"0B", x"5E", x"00", x"00", x"00", x"0B", x"68", x"00", x"00", x"00", x"0B", x"72", x"00", x"00", x"00", x"0B", x"7C", x"00", x"00", x"00", x"0B", x"86", x"00", x"00", x"00", x"0B", x"90", x"00", x"00", x"00", x"0B", x"9A", x"00", x"00", x"00", x"0B", x"A4", x"00", x"00", x"00", x"0B", x"AE", x"00", x"00", x"00", x"0B", x"B8", x"00", x"00", x"00", x"0B", x"C2", x"00", x"00", x"00", x"0B", x"CC", x"00", x"00", x"00", x"0B", x"D6", x"00", x"00", x"00", x"0B", x"E0", x"00", x"00", x"00", x"0B", x"EA", x"00", x"00", x"00", x"0B", x"F4", x"00", x"00", x"00", x"0B", x"FE", x"00", x"00", x"00", x"0C", x"08", x"00", x"00", x"00", x"0C", x"12", x"00", x"00", x"00", x"0C", x"1C", x"00", x"00", x"00", x"0C", x"26", x"00", x"00", x"00", x"0C", x"30", x"00", x"00", x"00", x"0C", x"3A", x"00", x"00", x"00", x"0C", x"44", x"00", x"00", x"00", x"0C", x"4E", x"00", x"00", x"00", x"0C", x"58", x"00", x"00", x"00", x"0C", x"62", x"00", x"00", x"00", x"0C", x"6C", x"00", x"00", x"00", x"0C", x"76", x"00", x"00", x"00", x"0C", x"80", x"00", x"00", x"00", x"0C", x"8A", x"00", x"00", x"00", x"0C", x"94", x"00", x"00", x"00", x"0C", x"9E", x"00", x"00", x"00", x"0C", x"A8", x"00", x"00", x"00", x"0C", x"B2", x"00", x"00", x"00", x"0C", x"BC", x"00", x"00", x"00", x"0C", x"C6", x"00", x"00", x"00", x"0C", x"D0", x"00", x"00", x"00", x"0C", x"DA", x"00", x"00", x"00", x"0C", x"E4", x"00", x"00", x"00", x"0C", x"EE", x"00", x"00", x"00", x"0C", x"F8", x"00", x"00", x"00", x"0D", x"02", x"00", x"00", x"00", x"0D", x"0C", x"00", x"00", x"00", x"0D", x"16", x"00", x"00", x"00", x"0D", x"20", x"00", x"00", x"00", x"0D", x"2A", x"00", x"00", x"00", x"0D", x"34", x"00", x"00", x"00", x"0D", x"3E", x"00", x"00", x"00", x"0D", x"48", x"00", x"00", x"00", x"0D", x"52", x"00", x"00", x"00", x"0D", x"5C", x"00", x"00", x"00", x"0D", x"66", x"00", x"00", x"00", x"0D", x"70", x"00", x"00", x"00", x"0D", x"7A", x"00", x"00", x"00", x"0D", x"84", x"00", x"00", x"00", x"0D", x"8E", x"00", x"00", x"00", x"0D", x"98", x"00", x"00", x"00", x"0D", x"A2", x"00", x"00", x"00", x"0D", x"AC", x"00", x"00", x"00", x"0D", x"B6", x"00", x"00", x"00", x"0D", x"C0", x"00", x"00", x"00", x"0D", x"CA", x"00", x"00", x"00", x"0D", x"D4", x"00", x"00", x"00", x"0D", x"DE", x"00", x"00", x"00", x"0D", x"E8", x"00", x"00", x"00", x"0D", x"F2", x"00", x"00", x"00", x"0D", x"FC", x"00", x"00", x"00", x"0E", x"06", x"00", x"00", x"00", x"0E", x"10", x"00", x"00", x"00", x"0E", x"1A", x"00", x"00", x"00", x"0E", x"24", x"00", x"00", x"00", x"0E", x"2E", x"00", x"00", x"00", x"0E", x"38", x"00", x"00", x"00", x"0E", x"42", x"00", x"00", x"00", x"0E", x"4C", x"00", x"00", x"00", x"0E", x"56", x"00", x"00", x"00", x"0E", x"60", x"00", x"00", x"00", x"0E", x"6A", x"00", x"00", x"00", x"0E", x"74", x"00", x"00", x"00", x"0E", x"7E", x"00", x"00", x"00", x"0E", x"88", x"00", x"00", x"00", x"0E", x"92", x"00", x"00", x"00", x"0E", x"9C", x"00", x"00", x"00", x"0E", x"A6", x"00", x"00", x"00", x"0E", x"B0", x"00", x"00", x"00", x"0E", x"BA", x"00", x"00", x"00", x"0E", x"C4", x"00", x"00", x"00", x"0E", x"CE", x"00", x"00", x"00", x"0E", x"D8", x"00", x"00", x"00", x"0E", x"E2", x"00", x"00", x"00", x"0E", x"EC", x"00", x"00", x"00", x"0E", x"F6", x"00", x"00", x"00", x"0F", x"00", x"00", x"00", x"00", x"0F", x"0A", x"00", x"00", x"00", x"0F", x"14", x"00", x"00", x"00", x"0F", x"1E", x"00", x"00", x"00", x"0F", x"28", x"00", x"00", x"00", x"0F", x"32", x"00", x"00", x"00", x"0F", x"3C", x"00", x"00", x"00", x"0F", x"46", x"00", x"00", x"00", x"0F", x"50", x"00", x"00", x"00", x"0F", x"5A", x"00", x"00", x"00", x"0F", x"64", x"00", x"00", x"00", x"0F", x"6E", x"00", x"00", x"00", x"0F", x"78", x"00", x"00", x"00", x"0F", x"82", x"00", x"00", x"00", x"0F", x"8C", x"00", x"00", x"00", x"0F", x"96", x"00", x"00", x"00", x"0F", x"A0", x"00", x"00", x"00", x"0F", x"AA", x"00", x"00", x"00", x"0F", x"B4", x"00", x"00", x"00", x"0F", x"BE", x"00", x"00", x"00", x"0F", x"C8", x"00", x"00", x"00", x"0F", x"D2", x"00", x"00", x"00", x"0F", x"DC", x"00", x"00", x"00", x"0F", x"E6", x"00", x"00", x"00", x"0F", x"F0", x"00", x"00", x"00", x"0F", x"FA", x"00", x"00", x"00", x"10", x"04", x"00", x"00", x"00", x"10", x"0E", x"00", x"00", x"00", x"10", x"18", x"00", x"00", x"00", x"10", x"22", x"00", x"00", x"00", x"10", x"2C", x"00", x"00", x"00", x"10", x"36", x"00", x"00", x"00", x"10", x"40", x"00", x"00", x"00", x"10", x"4A", x"00", x"00", x"00", x"10", x"54", x"00", x"00", x"00", x"10", x"5E", x"00", x"00", x"00", x"10", x"68", x"00", x"00", x"00", x"10", x"72", x"00", x"00", x"00", x"10", x"7C", x"00", x"00", x"00", x"10", x"86", x"00", x"00", x"00", x"10", x"90", x"00", x"00", x"00", x"10", x"9A", x"00", x"00", x"00", x"10", x"A4", x"00", x"00", x"00", x"10", x"AE", x"00", x"00", x"00", x"10", x"B8", x"00", x"00", x"00", x"10", x"C2", x"00", x"00", x"00", x"10", x"CC", x"00", x"00", x"00", x"10", x"D6", x"00", x"00", x"00", x"10", x"E0", x"00", x"00", x"00", x"10", x"EA", x"00", x"00", x"00", x"10", x"F4", x"00", x"00", x"00", x"10", x"FE", x"00", x"00", x"00", x"11", x"08", x"00", x"00", x"00", x"11", x"12", x"00", x"00", x"00", x"11", x"1C", x"00", x"00", x"00", x"11", x"26", x"00", x"00", x"00", x"11", x"30", x"00", x"00", x"00", x"11", x"3A", x"00", x"00", x"00", x"11", x"44", x"00", x"00", x"00", x"11", x"4E", x"00", x"00", x"00", x"11", x"58", x"00", x"00", x"00", x"11", x"62", x"00", x"00", x"00", x"11", x"6C", x"00", x"00", x"00", x"11", x"76", x"00", x"00", x"00", x"11", x"80", x"00", x"00", x"00", x"11", x"8A", x"00", x"00", x"00", x"11", x"94", x"00", x"00", x"00", x"11", x"9E", x"00", x"00", x"00", x"11", x"A8", x"00", x"00", x"00", x"11", x"B2", x"00", x"00", x"00", x"11", x"BC", x"00", x"00", x"00", x"11", x"C6", x"00", x"00", x"00", x"11", x"D0", x"00", x"00", x"00", x"11", x"DA", x"00", x"00", x"00", x"11", x"E4", x"00", x"00", x"00", x"11", x"EE", x"00", x"00", x"00", x"11", x"F8", x"00", x"00", x"00", x"12", x"02", x"00", x"00", x"00", x"12", x"0C", x"00", x"00", x"00", x"12", x"16", x"00", x"00", x"00", x"12", x"20", x"00", x"00", x"00", x"12", x"2A", x"00", x"00", x"00", x"12", x"34", x"00", x"00", x"00", x"12", x"3E", x"00", x"00", x"00", x"12", x"48", x"00", x"00", x"00", x"12", x"52", x"00", x"00", x"00", x"12", x"5C", x"00", x"00", x"00", x"12", x"66", x"00", x"00", x"00", x"12", x"70", x"00", x"00", x"00", x"12", x"7A", x"00", x"00", x"00", x"12", x"84", x"00", x"00", x"00", x"12", x"8E", x"00", x"00", x"00", x"12", x"98", x"00", x"00", x"00", x"12", x"A2", x"00", x"00", x"00", x"12", x"AC", x"00", x"00", x"00", x"12", x"B6", x"00", x"00", x"00", x"12", x"C0", x"00", x"00", x"00", x"12", x"CA", x"00", x"00", x"00", x"12", x"D4", x"00", x"00", x"00", x"12", x"DE", x"00", x"00", x"00", x"12", x"E8", x"00", x"00", x"00", x"12", x"F2", x"00", x"00", x"00", x"12", x"FC", x"00", x"00", x"00", x"13", x"06", x"00", x"00", x"00", x"13", x"10", x"00", x"00", x"00", x"13", x"1A", x"00", x"00", x"00", x"13", x"24", x"00", x"00", x"00", x"13", x"2E", x"00", x"00", x"00", x"13", x"38", x"00", x"00", x"00", x"13", x"42", x"00", x"00", x"00", x"13", x"4C", x"00", x"00", x"00", x"13", x"56", x"00", x"00", x"00", x"13", x"60", x"00", x"00", x"00", x"13", x"6A", x"00", x"00", x"00", x"13", x"74", x"00", x"00", x"00", x"13", x"7E", x"00", x"00", x"00", x"13", x"88", x"00", x"00", x"00", x"13", x"92", x"00", x"00", x"00", x"13", x"9C", x"00", x"00", x"00", x"13", x"A6", x"00", x"00", x"00", x"13", x"B0", x"00", x"00", x"00", x"13", x"BA", x"00", x"00", x"00", x"13", x"C4", x"00", x"00", x"00", x"13", x"CE", x"00", x"00", x"00", x"13", x"D8", x"00", x"00", x"00", x"13", x"E2", x"00", x"00", x"00", x"13", x"EC", x"00", x"00", x"00", x"13", x"F6", x"00", x"00", x"00", x"14", x"00", x"00", x"00", x"00", x"14", x"0A", x"00", x"00", x"00", x"14", x"14", x"00", x"00", x"00", x"14", x"1E", x"00", x"00", x"00", x"14", x"28", x"00", x"00", x"00", x"14", x"32", x"00", x"00", x"00", x"14", x"3C", x"00", x"00", x"00", x"14", x"46", x"00", x"00", x"00", x"14", x"50", x"00", x"00", x"00", x"14", x"5A", x"00", x"00", x"00", x"14", x"64", x"00", x"00", x"00", x"14", x"6E", x"00", x"00", x"00", x"14", x"78", x"00", x"00", x"00", x"14", x"82", x"00", x"00", x"00", x"14", x"8C", x"00", x"00", x"00", x"14", x"96", x"00", x"00", x"00", x"14", x"A0", x"00", x"00", x"00", x"14", x"AA", x"00", x"00", x"00", x"14", x"B4", x"00", x"00", x"00", x"14", x"BE", x"00", x"00", x"00", x"14", x"C8", x"00", x"00", x"00", x"14", x"D2", x"00", x"00", x"00", x"14", x"DC", x"00", x"00", x"00", x"14", x"E6", x"00", x"00", x"00", x"14", x"F0", x"00", x"00", x"00", x"14", x"FA", x"00", x"00", x"00", x"15", x"04", x"00", x"00", x"00", x"15", x"0E", x"00", x"00", x"00", x"15", x"18", x"00", x"00", x"00", x"15", x"22", x"00", x"00", x"00", x"15", x"2C", x"00", x"00", x"00", x"15", x"36", x"00", x"00", x"00", x"15", x"40", x"00", x"00", x"00", x"15", x"4A", x"00", x"00", x"00", x"15", x"54", x"00", x"00", x"00", x"15", x"5E", x"00", x"00", x"00", x"15", x"68", x"00", x"00", x"00", x"15", x"72", x"00", x"00", x"00", x"15", x"7C", x"00", x"00", x"00", x"15", x"86", x"00", x"00", x"00", x"15", x"90", x"00", x"00", x"00", x"15", x"9A", x"00", x"00", x"00", x"15", x"A4", x"00", x"00", x"00", x"15", x"AE", x"00", x"00", x"00", x"15", x"B8", x"00", x"00", x"00", x"15", x"C2", x"00", x"00", x"00", x"15", x"CC", x"00", x"00", x"00", x"15", x"D6", x"00", x"00", x"00", x"15", x"E0", x"00", x"00", x"00", x"15", x"EA", x"00", x"00", x"00", x"15", x"F4", x"00", x"00", x"00", x"15", x"FE", x"00", x"00", x"00", x"16", x"08", x"00", x"00", x"00", x"16", x"12", x"00", x"00", x"00", x"16", x"1C", x"00", x"00", x"00", x"16", x"26", x"00", x"00", x"00", x"16", x"30", x"00", x"00", x"00", x"16", x"3A", x"00", x"00", x"00", x"16", x"44", x"00", x"00", x"00", x"16", x"4E", x"00", x"00", x"00", x"16", x"58", x"00", x"00", x"00", x"16", x"62", x"00", x"00", x"00", x"16", x"6C", x"00", x"00", x"00", x"16", x"76", x"00", x"00", x"00", x"16", x"80", x"00", x"00", x"00", x"16", x"8A", x"00", x"00", x"00", x"16", x"94", x"00", x"00", x"00", x"16", x"9E", x"00", x"00", x"00", x"16", x"A8", x"00", x"00", x"00", x"16", x"B2", x"00", x"00", x"00", x"16", x"BC", x"00", x"00", x"00", x"16", x"C6", x"00", x"00", x"00", x"16", x"D0", x"00", x"00", x"00", x"16", x"DA", x"00", x"00", x"00", x"16", x"E4", x"00", x"00", x"00", x"16", x"EE", x"00", x"00", x"00", x"16", x"F8", x"00", x"00", x"00", x"17", x"02", x"00", x"00", x"00", x"17", x"0C", x"00", x"00", x"00", x"17", x"16", x"00", x"00", x"00", x"17", x"20", x"00", x"00", x"00", x"17", x"2A", x"00", x"00", x"00", x"17", x"34", x"00", x"00", x"00", x"17", x"3E", x"00", x"00", x"00", x"17", x"48", x"00", x"00", x"00", x"17", x"52", x"00", x"00", x"00", x"17", x"5C", x"00", x"00", x"00", x"17", x"66", x"00", x"00", x"00", x"17", x"70", x"00", x"00", x"00", x"17", x"7A", x"00", x"00", x"00", x"17", x"84", x"00", x"00", x"00", x"17", x"8E", x"00", x"00", x"00", x"17", x"98", x"00", x"00", x"00", x"17", x"A2", x"00", x"00", x"00", x"17", x"AC", x"00", x"00", x"00", x"17", x"B6", x"00", x"00", x"00", x"17", x"C0", x"00", x"00", x"00", x"17", x"CA", x"00", x"00", x"00", x"17", x"D4", x"00", x"00", x"00", x"17", x"DE", x"00", x"00", x"00", x"17", x"E8", x"00", x"00", x"00", x"17", x"F2", x"00", x"00", x"00", x"17", x"FC", x"00", x"00", x"00", x"18", x"06", x"00", x"00", x"00", x"18", x"10", x"00", x"00", x"00", x"18", x"1A", x"00", x"00", x"00", x"18", x"24", x"00", x"00", x"00", x"18", x"2E", x"00", x"00", x"00", x"18", x"38", x"00", x"00", x"00", x"18", x"42", x"00", x"00", x"00", x"18", x"4C", x"00", x"00", x"00", x"18", x"56", x"00", x"00", x"00", x"18", x"60", x"00", x"00", x"00", x"18", x"6A", x"00", x"00", x"00", x"18", x"74", x"00", x"00", x"00", x"18", x"7E", x"00", x"00", x"00", x"18", x"88", x"00", x"00", x"00", x"18", x"92", x"00", x"00", x"00", x"18", x"9C", x"00", x"00", x"00", x"18", x"A6", x"00", x"00", x"00", x"18", x"B0", x"00", x"00", x"00", x"18", x"BA", x"00", x"00", x"00", x"18", x"C4", x"00", x"00", x"00", x"18", x"CE", x"00", x"00", x"00", x"18", x"D8", x"00", x"00", x"00", x"18", x"E2", x"00", x"00", x"00", x"18", x"EC", x"00", x"00", x"00", x"18", x"F6", x"00", x"00", x"00", x"19", x"00", x"00", x"00", x"00", x"19", x"0A", x"00", x"00", x"00", x"19", x"14", x"00", x"00", x"00", x"19", x"1E", x"00", x"00", x"00", x"19", x"28", x"00", x"00", x"00", x"19", x"32", x"00", x"00", x"00", x"19", x"3C", x"00", x"00", x"00", x"19", x"46", x"00", x"00", x"00", x"19", x"50", x"00", x"00", x"00", x"19", x"5A", x"00", x"00", x"00", x"19", x"64", x"00", x"00", x"00", x"19", x"6E", x"00", x"00", x"00", x"19", x"78", x"00", x"00", x"00", x"19", x"82", x"00", x"00", x"00", x"19", x"8C", x"00", x"00", x"00", x"19", x"96", x"00", x"00", x"00", x"19", x"A0", x"00", x"00", x"00", x"19", x"AA", x"00", x"00", x"00", x"19", x"B4", x"00", x"00", x"00", x"19", x"BE", x"00", x"00", x"00", x"19", x"C8", x"00", x"00", x"00", x"19", x"D2", x"00", x"00", x"00", x"19", x"DC", x"00", x"00", x"00", x"19", x"E6", x"00", x"00", x"00", x"19", x"F0", x"00", x"00", x"00", x"19", x"FA", x"00", x"00", x"00", x"1A", x"04", x"00", x"00", x"00", x"1A", x"0E", x"00", x"00", x"00", x"1A", x"18", x"00", x"00", x"00", x"1A", x"22", x"00", x"00", x"00", x"1A", x"2C", x"00", x"00", x"00", x"1A", x"36", x"00", x"00", x"00", x"1A", x"40", x"00", x"00", x"00", x"1A", x"4A", x"00", x"00", x"00", x"1A", x"54", x"00", x"00", x"00", x"1A", x"5E", x"00", x"00", x"00", x"1A", x"68", x"00", x"00", x"00", x"1A", x"72", x"00", x"00", x"00", x"1A", x"7C", x"00", x"00", x"00", x"1A", x"86", x"00", x"00", x"00", x"1A", x"90", x"00", x"00", x"00", x"1A", x"9A", x"00", x"00", x"00", x"1A", x"A4", x"00", x"00", x"00", x"1A", x"AE", x"00", x"00", x"00", x"1A", x"B8", x"00", x"00", x"00", x"1A", x"C2", x"00", x"00", x"00", x"1A", x"CC", x"00", x"00", x"00", x"1A", x"D6", x"00", x"00", x"00", x"1A", x"E0", x"00", x"00", x"00", x"1A", x"EA", x"00", x"00", x"00", x"1A", x"F4", x"00", x"00", x"00", x"1A", x"FE", x"00", x"00", x"00", x"1B", x"08", x"00", x"00", x"00", x"1B", x"12", x"00", x"00", x"00", x"1B", x"1C", x"00", x"00", x"00", x"1B", x"26", x"00", x"00", x"00", x"1B", x"30", x"00", x"00", x"00", x"1B", x"3A", x"00", x"00", x"00", x"1B", x"44", x"00", x"00", x"00", x"1B", x"4E", x"00", x"00", x"00", x"1B", x"58", x"00", x"00", x"00", x"1B", x"62", x"00", x"00", x"00", x"1B", x"6C", x"00", x"00", x"00", x"1B", x"76", x"00", x"00", x"00", x"1B", x"80", x"00", x"00", x"00", x"1B", x"8A", x"00", x"00", x"00", x"1B", x"94", x"00", x"00", x"00", x"1B", x"9E", x"00", x"00", x"00", x"1B", x"A8", x"00", x"00", x"00", x"1B", x"B2", x"00", x"00", x"00", x"1B", x"BC", x"00", x"00", x"00", x"1B", x"C6", x"00", x"00", x"00", x"1B", x"D0", x"00", x"00", x"00", x"1B", x"DA", x"00", x"00", x"00", x"1B", x"E4", x"00", x"00", x"00", x"1B", x"EE", x"00", x"00", x"00", x"1B", x"F8", x"00", x"00", x"00", x"1C", x"02", x"00", x"00", x"00", x"1C", x"0C", x"00", x"00", x"00", x"1C", x"16", x"00", x"00", x"00", x"1C", x"20", x"00", x"00", x"00", x"1C", x"2A", x"00", x"00", x"00", x"1C", x"34", x"00", x"00", x"00", x"1C", x"3E", x"00", x"00", x"00", x"1C", x"48", x"00", x"00", x"00", x"1C", x"52", x"00", x"00", x"00", x"1C", x"5C", x"00", x"00", x"00", x"1C", x"66", x"00", x"00", x"00", x"1C", x"70", x"00", x"00", x"00", x"1C", x"7A", x"00", x"00", x"00", x"1C", x"84", x"00", x"00", x"00", x"1C", x"8E", x"00", x"00", x"00", x"1C", x"98", x"00", x"00", x"00", x"1C", x"A2", x"00", x"00", x"00", x"1C", x"AC", x"00", x"00", x"00", x"1C", x"B6", x"00", x"00", x"00", x"1C", x"C0", x"00", x"00", x"00", x"1C", x"CA", x"00", x"00", x"00", x"1C", x"D4", x"00", x"00", x"00", x"1C", x"DE", x"00", x"00", x"00", x"1C", x"E8", x"00", x"00", x"00", x"1C", x"F2", x"00", x"00", x"00", x"1C", x"FC", x"00", x"00", x"00", x"1D", x"06", x"00", x"00", x"00", x"1D", x"10", x"00", x"00", x"00", x"1D", x"1A", x"00", x"00", x"00", x"1D", x"24", x"00", x"00", x"00", x"1D", x"2E", x"00", x"00", x"00", x"1D", x"38", x"00", x"00", x"00", x"1D", x"42", x"00", x"00", x"00", x"1D", x"4C", x"00", x"00", x"00", x"1D", x"56", x"00", x"00", x"00", x"1D", x"60", x"00", x"00", x"00", x"1D", x"6A", x"00", x"00", x"00", x"1D", x"74", x"00", x"00", x"00", x"1D", x"7E", x"00", x"00", x"00", x"1D", x"88", x"00", x"00", x"00", x"1D", x"92", x"00", x"00", x"00", x"1D", x"9C", x"00", x"00", x"00", x"1D", x"A6", x"00", x"00", x"00", x"1D", x"B0", x"00", x"00", x"00", x"1D", x"BA", x"00", x"00", x"00", x"1D", x"C4", x"00", x"00", x"00", x"1D", x"CE", x"00", x"00", x"00", x"1D", x"D8", x"00", x"00", x"00", x"1D", x"E2", x"00", x"00", x"00", x"1D", x"EC", x"00", x"00", x"00", x"1D", x"F6", x"00", x"00", x"00", x"1E", x"00", x"00", x"00", x"00", x"1E", x"0A", x"00", x"00", x"00", x"1E", x"14", x"00", x"00", x"00", x"1E", x"1E", x"00", x"00", x"00", x"1E", x"28", x"00", x"00", x"00", x"1E", x"32", x"00", x"00", x"00", x"1E", x"3C", x"00", x"00", x"00", x"1E", x"46", x"00", x"00", x"00", x"1E", x"50", x"00", x"00", x"00", x"1E", x"5A", x"00", x"00", x"00", x"1E", x"64", x"00", x"00", x"00", x"1E", x"6E", x"00", x"00", x"00", x"1E", x"78", x"00", x"00", x"00", x"1E", x"82", x"00", x"00", x"00", x"1E", x"8C", x"00", x"00", x"00", x"1E", x"96", x"00", x"00", x"00", x"1E", x"A0", x"00", x"00", x"00", x"1E", x"AA", x"00", x"00", x"00", x"1E", x"B4", x"00", x"00", x"00", x"1E", x"BE", x"00", x"00", x"00", x"1E", x"C8", x"00", x"00", x"00", x"1E", x"D2", x"00", x"00", x"00", x"1E", x"DC", x"00", x"00", x"00", x"1E", x"E6", x"00", x"00", x"00", x"1E", x"F0", x"00", x"00", x"00", x"1E", x"FA", x"00", x"00", x"00", x"1F", x"04", x"00", x"00", x"00", x"1F", x"0E", x"00", x"00", x"00", x"1F", x"18", x"00", x"00", x"00", x"1F", x"22", x"00", x"00", x"00", x"1F", x"2C", x"00", x"00", x"00", x"1F", x"36", x"00", x"00", x"00", x"1F", x"40", x"00", x"00", x"00", x"1F", x"4A", x"00", x"00", x"00", x"1F", x"54", x"00", x"00", x"00", x"1F", x"5E", x"00", x"00", x"00", x"1F", x"68", x"00", x"00", x"00", x"1F", x"72", x"00", x"00", x"00", x"1F", x"7C", x"00", x"00", x"00", x"1F", x"86", x"00", x"00", x"00", x"1F", x"90", x"00", x"00", x"00", x"1F", x"9A", x"00", x"00", x"00", x"1F", x"A4", x"00", x"00", x"00", x"1F", x"AE", x"00", x"00", x"00", x"1F", x"B8", x"00", x"00", x"00", x"1F", x"C2", x"00", x"00", x"00", x"1F", x"CC", x"00", x"00", x"00", x"1F", x"D6", x"00", x"00", x"00", x"1F", x"E0", x"00", x"00", x"00", x"1F", x"EA", x"00", x"00", x"00", x"1F", x"F4", x"00", x"00", x"00", x"1F", x"FE", x"00", x"00", x"00", x"20", x"08", x"00", x"00", x"00", x"20", x"12", x"00", x"00", x"00", x"20", x"1C", x"00", x"00", x"00", x"20", x"26", x"00", x"00", x"00", x"20", x"30", x"00", x"00", x"00", x"20", x"3A", x"00", x"00", x"00", x"20", x"44", x"00", x"00", x"00", x"20", x"4E", x"00", x"00", x"00", x"20", x"58", x"00", x"00", x"00", x"20", x"62", x"00", x"00", x"00", x"20", x"6C", x"00", x"00", x"00", x"20", x"76", x"00", x"00", x"00", x"20", x"80", x"00", x"00", x"00", x"20", x"8A", x"00", x"00", x"00", x"20", x"94", x"00", x"00", x"00", x"20", x"9E", x"00", x"00", x"00", x"20", x"A8", x"00", x"00", x"00", x"20", x"B2", x"00", x"00", x"00", x"20", x"BC", x"00", x"00", x"00", x"20", x"C6", x"00", x"00", x"00", x"20", x"D0", x"00", x"00", x"00", x"20", x"DA", x"00", x"00", x"00", x"20", x"E4", x"00", x"00", x"00", x"20", x"EE", x"00", x"00", x"00", x"20", x"F8", x"00", x"00", x"00", x"21", x"02", x"00", x"00", x"00", x"21", x"0C", x"00", x"00", x"00", x"21", x"16", x"00", x"00", x"00", x"21", x"20", x"00", x"00", x"00", x"21", x"2A", x"00", x"00", x"00", x"21", x"34", x"00", x"00", x"00", x"21", x"3E", x"00", x"00", x"00", x"21", x"48", x"00", x"00", x"00", x"21", x"52", x"00", x"00", x"00", x"21", x"5C", x"00", x"00", x"00", x"21", x"66", x"00", x"00", x"00", x"21", x"70", x"00", x"00", x"00", x"21", x"7A", x"00", x"00", x"00", x"21", x"84", x"00", x"00", x"00", x"21", x"8E", x"00", x"00", x"00", x"21", x"98", x"00", x"00", x"00", x"21", x"A2", x"00", x"00", x"00", x"21", x"AC", x"00", x"00", x"00", x"21", x"B6", x"00", x"00", x"00", x"21", x"C0", x"00", x"00", x"00", x"21", x"CA", x"00", x"00", x"00", x"21", x"D4", x"00", x"00", x"00", x"21", x"DE", x"00", x"00", x"00", x"21", x"E8", x"00", x"00", x"00", x"21", x"F2", x"00", x"00", x"00", x"21", x"FC", x"00", x"00", x"00", x"22", x"06", x"00", x"00", x"00", x"22", x"10", x"00", x"00", x"00", x"22", x"1A", x"00", x"00", x"00", x"22", x"24", x"00", x"00", x"00", x"22", x"2E", x"00", x"00", x"00", x"22", x"38", x"00", x"00", x"00", x"22", x"42", x"00", x"00", x"00", x"22", x"4C", x"00", x"00", x"00", x"22", x"56", x"00", x"00", x"00", x"22", x"60", x"00", x"00", x"00", x"22", x"6A", x"00", x"00", x"00", x"22", x"74", x"00", x"00", x"00", x"22", x"7E", x"00", x"00", x"00", x"22", x"88", x"00", x"00", x"00", x"22", x"92", x"00", x"00", x"00", x"22", x"9C", x"00", x"00", x"00", x"22", x"A6", x"00", x"00", x"00", x"22", x"B0", x"00", x"00", x"00", x"22", x"BA", x"00", x"00", x"00", x"22", x"C4", x"00", x"00", x"00", x"22", x"CE", x"00", x"00", x"00", x"22", x"D8", x"00", x"00", x"00", x"22", x"E2", x"00", x"00", x"00", x"22", x"EC", x"00", x"00", x"00", x"22", x"F6", x"00", x"00", x"00", x"23", x"00", x"00", x"00", x"00", x"23", x"0A", x"00", x"00", x"00", x"23", x"14", x"00", x"00", x"00", x"23", x"1E", x"00", x"00", x"00", x"23", x"28", x"00", x"00", x"00", x"23", x"32", x"00", x"00", x"00", x"23", x"3C", x"00", x"00", x"00", x"23", x"46", x"00", x"00", x"00", x"23", x"50", x"00", x"00", x"00", x"23", x"5A", x"00", x"00", x"00", x"23", x"64", x"00", x"00", x"00", x"23", x"6E", x"00", x"00", x"00", x"23", x"78", x"00", x"00", x"00", x"23", x"82", x"00", x"00", x"00", x"23", x"8C", x"00", x"00", x"00", x"23", x"96", x"00", x"00", x"00", x"23", x"A0", x"00", x"00", x"00", x"23", x"AA", x"00", x"00", x"00", x"23", x"B4", x"00", x"00", x"00", x"23", x"BE", x"00", x"00", x"00", x"23", x"C8", x"00", x"00", x"00", x"23", x"D2", x"00", x"00", x"00", x"23", x"DC", x"00", x"00", x"00", x"23", x"E6", x"00", x"00", x"00", x"23", x"F0", x"00", x"00", x"00", x"23", x"FA", x"00", x"00", x"00", x"24", x"04", x"00", x"00", x"00", x"24", x"0E", x"00", x"00", x"00", x"24", x"18", x"00", x"00", x"00", x"24", x"22", x"00", x"00", x"00", x"24", x"2C", x"00", x"00", x"00", x"24", x"36", x"00", x"00", x"00", x"24", x"40", x"00", x"00", x"00", x"24", x"4A", x"00", x"00", x"00", x"24", x"54", x"00", x"00", x"00", x"24", x"5E", x"00", x"00", x"00", x"24", x"68", x"00", x"00", x"00", x"24", x"72", x"00", x"00", x"00", x"24", x"7C", x"00", x"00", x"00", x"24", x"86", x"00", x"00", x"00", x"24", x"90", x"00", x"00", x"00", x"24", x"9A", x"00", x"00", x"00", x"24", x"A4", x"00", x"00", x"00", x"24", x"AE", x"00", x"00", x"00", x"24", x"B8", x"00", x"00", x"00", x"24", x"C2", x"00", x"00", x"00", x"24", x"CC", x"00", x"00", x"00", x"24", x"D6", x"00", x"00", x"00", x"24", x"E0", x"00", x"00", x"00", x"24", x"EA", x"00", x"00", x"00", x"24", x"F4", x"00", x"00", x"00", x"24", x"FE", x"00", x"00", x"00", x"25", x"08", x"00", x"00", x"00", x"25", x"12", x"00", x"00", x"00", x"25", x"1C", x"00", x"00", x"00", x"25", x"26", x"00", x"00", x"00", x"25", x"30", x"00", x"00", x"00", x"25", x"3A", x"00", x"00", x"00", x"25", x"44", x"00", x"00", x"00", x"25", x"4E", x"00", x"00", x"00", x"25", x"58", x"00", x"00", x"00", x"25", x"62", x"00", x"00", x"00", x"25", x"6C", x"00", x"00", x"00", x"25", x"76", x"00", x"00", x"00", x"25", x"80", x"00", x"00", x"00", x"25", x"8A", x"00", x"00", x"00", x"25", x"94", x"00", x"00", x"00", x"25", x"9E", x"00", x"00", x"00", x"25", x"A8", x"00", x"00", x"00", x"25", x"B2", x"00", x"00", x"00", x"25", x"BC", x"00", x"00", x"00", x"25", x"C6", x"00", x"00", x"00", x"25", x"D0", x"00", x"00", x"00", x"25", x"DA", x"00", x"00", x"00", x"25", x"E4", x"00", x"00", x"00", x"25", x"EE", x"00", x"00", x"00", x"25", x"F8", x"00", x"00", x"00", x"26", x"02", x"00", x"00", x"00", x"26", x"0C", x"00", x"00", x"00", x"26", x"16", x"00", x"00", x"00", x"26", x"20", x"00", x"00", x"00", x"26", x"2A", x"00", x"00", x"00", x"26", x"34", x"00", x"00", x"00", x"26", x"3E", x"00", x"00", x"00", x"26", x"48", x"00", x"00", x"00", x"26", x"52", x"00", x"00", x"00", x"26", x"5C", x"00", x"00", x"00", x"26", x"66", x"00", x"00", x"00", x"26", x"70", x"00", x"00", x"00", x"26", x"7A", x"00", x"00", x"00", x"26", x"84", x"00", x"00", x"00", x"26", x"8E", x"00", x"00", x"00", x"26", x"98", x"00", x"00", x"00", x"26", x"A2", x"00", x"00", x"00", x"26", x"AC", x"00", x"00", x"00", x"26", x"B6", x"00", x"00", x"00", x"26", x"C0", x"00", x"00", x"00", x"26", x"CA", x"00", x"00", x"00", x"26", x"D4", x"00", x"00", x"00", x"26", x"DE", x"00", x"00", x"00", x"26", x"E8", x"00", x"00", x"00", x"26", x"F2", x"00", x"00", x"00", x"26", x"FC", x"00", x"00", x"00", x"27", x"06", x"00", x"00", x"00", x"27", x"10", x"00", x"00", x"00", x"27", x"1A", x"00", x"00", x"00", x"27", x"24", x"00", x"00", x"00", x"27", x"2E", x"00", x"00", x"00", x"27", x"38", x"00", x"00", x"00", x"27", x"42", x"00", x"00", x"00", x"27", x"4C", x"00", x"00", x"00", x"27", x"56", x"00", x"00", x"00", x"27", x"60", x"00", x"00", x"00", x"27", x"6A", x"00", x"00", x"00", x"27", x"74", x"00", x"00", x"00", x"27", x"7E", x"00", x"00", x"00", x"27", x"88", x"00", x"00", x"00", x"27", x"92", x"00", x"00", x"00", x"27", x"9C", x"00", x"00", x"00", x"27", x"A6", x"00", x"00", x"00", x"27", x"B0", x"00", x"00", x"00", x"27", x"BA", x"00", x"00", x"00", x"27", x"C4", x"00", x"00", x"00", x"27", x"CE", x"00", x"00", x"00", x"27", x"D8", x"00", x"00", x"00", x"27", x"E2", x"00", x"00", x"00", x"27", x"EC", x"00", x"00", x"00", x"27", x"F6", x"00", x"00");

type Tseq_array3 is array (0 to 42+5-1) of std_logic_vector(7 downto 0);
constant seq_array3:Tseq_array3:=(x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"16", x"ea", x"ca", x"09", x"3a", x"08", x"00", x"45", x"00", x"00", x"1f", x"57", x"ac", x"00", x"00", x"80", x"11", x"21", x"74", x"c0", x"a8", x"01", x"06", x"ff", x"ff", x"ff", x"ff", x"e2", x"ce", x"ec", x"be", x"00", x"0b", x"14", x"9c",
x"A5", x"04", x"02", x"00", x"30");

type Tseq_array4 is array (0 to 42+16-1) of std_logic_vector(7 downto 0);
constant seq_array4:Tseq_array4:=(x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"00", x"16", x"ea", x"ca", x"09", x"3a", x"08", x"00", x"45", x"00", x"00", x"1f", x"57", x"ac", x"00", x"00", x"80", x"11", x"21", x"74", x"c0", x"a8", x"01", x"06", x"ff", x"ff", x"ff", x"ff", x"e2", x"ce", x"ec", x"be", x"00", x"0b", x"14", x"9c",
x"A5", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");

constant RESP_NUM:natural:=5;
type Tsizes is array(0 to 5-1) of integer;
constant sizes:Tsizes:=(58, 47, 10290, 47, 58);
type Tstm is (FINISH,TX_STATE0, TX_STATE1, TX_STATE2, TX_STATE3, TX_STATE4,WAIT_RESPONSE0, WAIT_RESPONSE1, WAIT_RESPONSE2, WAIT_RESPONSE3, WAIT_RESPONSE4,START_DELAY0, START_DELAY1, START_DELAY2, START_DELAY3, START_DELAY4);
signal stm:Tstm;

begin

process(clk)
begin
	if rising_edge(clk) then
		if reset='1' then
			stm<=WAIT_RESPONSE0;
			delay_cnt<=(others=>'1');
			dv_o<='0';
		elsif ce='1' then    --# reset
			case stm is
			when WAIT_RESPONSE0=>
				if can_go='1' then
					stm<=START_DELAY0;
				end if;
				delay_cnt<=(others=>'1');
				dv_o<='0';
			when START_DELAY0=>	
				if unsigned(delay_cnt)>0 then
					delay_cnt<=delay_cnt-1;
				else
					stm<=TX_STATE0;
				end if;
				cnt<=0;
				dv_o<='0';
			when TX_STATE0=>
				dv_o<='1';
				data_o<=seq_array0(cnt);
					if cnt<sizes(0)-1 then
						cnt<=cnt+1;
					else
						stm<=WAIT_RESPONSE1;
					end if;
			when WAIT_RESPONSE1=>
				if can_go='1' then
					stm<=START_DELAY1;
				end if;
				delay_cnt<=(others=>'1');
				dv_o<='0';
			when START_DELAY1=>	
				if unsigned(delay_cnt)>0 then
					delay_cnt<=delay_cnt-1;
				else
					stm<=TX_STATE1;
				end if;
				cnt<=0;
				dv_o<='0';
			when TX_STATE1=>
				dv_o<='1';
				data_o<=seq_array1(cnt);
					if cnt<sizes(1)-1 then
						cnt<=cnt+1;
					else
						stm<=WAIT_RESPONSE2;
					end if;
			when WAIT_RESPONSE2=>
				if can_go='1' then
					stm<=START_DELAY2;
				end if;
				delay_cnt<=(others=>'1');
				dv_o<='0';
			when START_DELAY2=>	
				if unsigned(delay_cnt)>0 then
					delay_cnt<=delay_cnt-1;
				else
					stm<=TX_STATE2;
				end if;
				cnt<=0;
				dv_o<='0';
			when TX_STATE2=>
				dv_o<='1';
				data_o<=seq_array2(cnt);
					if cnt<sizes(2)-1 then
						cnt<=cnt+1;
					else
						stm<=WAIT_RESPONSE3;
					end if;
			when WAIT_RESPONSE3=>
				if can_go='1' then
					stm<=START_DELAY3;
				end if;
				delay_cnt<=(others=>'1');
				dv_o<='0';
			when START_DELAY3=>	
				if unsigned(delay_cnt)>0 then
					delay_cnt<=delay_cnt-1;
				else
					stm<=TX_STATE3;
				end if;
				cnt<=0;
				dv_o<='0';
			when TX_STATE3=>
				dv_o<='1';
				data_o<=seq_array3(cnt);
					if cnt<sizes(3)-1 then
						cnt<=cnt+1;
					else
						stm<=WAIT_RESPONSE4;
					end if;
			when WAIT_RESPONSE4=>
				if can_go='1' then
					stm<=START_DELAY4;
				end if;
				delay_cnt<=(others=>'1');
				dv_o<='0';
			when START_DELAY4=>	
				if unsigned(delay_cnt)>0 then
					delay_cnt<=delay_cnt-1;
				else
					stm<=TX_STATE4;
				end if;
				cnt<=0;
				dv_o<='0';
			when TX_STATE4=>
				dv_o<='1';
				data_o<=seq_array4(cnt);
					if cnt<sizes(4)-1 then
						cnt<=cnt+1;
					else
					stm<=FINISH;
					end if;
			when FINISH=>
				 dv_o<='0';
				 data_o<=x"00";
			when others=>
			end case;
		end if; --# reset
	end if;
end process;

end cpp_response2vhdl;
