---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
--  version		: $Version:	1.0 $ 
--  revision		: $Revision: 1.1.1.1 $ 
--  designer name  	: $Author: jzhang $ 
--  company name   	: altera corp.
--  company address	: 101 innovation drive
--                  	  san jose, california 95134
--                  	  u.s.a.
-- 
--  copyright altera corp. 2003
-- 
-- 
--  $Header: /ipbu/cvs/dsp/projects/FFT/src/rtl/lib/asj_fft_mult_add.vhd,v 1.1.1.1 2005/12/08 01:14:15 jzhang Exp $ 
--  $log$ 
--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------- 
-- megafunction wizard: %ALTMULT_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTMULT_ADD 

-- ============================================================
-- File Name: asj_fft_cmults_std.vhd
-- Megafunction Name(s):
-- 			ALTMULT_ADD
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
-- ************************************************************


--Copyright (C) 1991-2003 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all; 

library work;
use work.fft_pack.all;
library lpm;
use lpm.lpm_components.all;
library altera_mf;
use altera_mf.altera_mf_components.all;


entity asj_fft_mult_add is
	generic(
		mpr : integer :=16;
		twr : integer :=12;
		dirn : string :="SUB"
	);
	port
	(
		clock0		: in std_logic  := '1';
		dataa_0		: in std_logic_vector (mpr-1 downto 0);
		dataa_1		: in std_logic_vector (mpr-1 downto 0);
		datab_0		: in std_logic_vector (twr-1 downto 0);
		datab_1		: in std_logic_vector (twr-1 downto 0);
		result		: out std_logic_vector (twr+mpr downto 0)
	);
end asj_fft_mult_add;


architecture syn of asj_fft_mult_add is
	
	ATTRIBUTE ALTERA_INTERNAL_OPTION : string;
	ATTRIBUTE ALTERA_INTERNAL_OPTION OF SYN : ARCHITECTURE IS "DSP_BLOCK_BALANCING=OFF";

	signal sub_wire0	: std_logic_vector (twr+mpr downto 0);
	signal sub_wire1	: std_logic_vector (mpr-1 downto 0);
	signal sub_wire2	: std_logic_vector (2*mpr-1 downto 0);
	signal sub_wire3	: std_logic_vector (mpr-1 downto 0);
	signal sub_wire4	: std_logic_vector (twr-1 downto 0);
	signal sub_wire5	: std_logic_vector (2*twr-1 downto 0);
	signal sub_wire6	: std_logic_vector (twr-1 downto 0);



	COMPONENT altmult_add
	GENERIC (
		input_register_a1		: STRING;
		multiplier_register0		: STRING;
		signed_pipeline_aclr_b		: STRING;
		multiplier_register1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		signed_aclr_a		: STRING;
		signed_register_a		: STRING;
		number_of_multipliers		: NATURAL;
		multiplier_aclr0		: STRING;
		signed_aclr_b		: STRING;
		signed_register_b		: STRING;
		lpm_type		: STRING;
		multiplier_aclr1		: STRING;
		input_aclr_b0		: STRING;
		output_register		: STRING;
		representation_a		: STRING;
		signed_pipeline_register_a		: STRING;
		width_result		: NATURAL;
		input_source_b0		: STRING;
		input_aclr_b1		: STRING;
		input_aclr_a0		: STRING;
		addnsub_multiplier_register1		: STRING;
		representation_b		: STRING;
		signed_pipeline_register_b		: STRING;
		input_source_b1		: STRING;
		input_source_a0		: STRING;
		input_aclr_a1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_source_a1		: STRING;
		addnsub_multiplier_aclr1		: STRING;
		output_aclr		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		width_a		: NATURAL;
		input_register_b0		: STRING;
		width_b		: NATURAL;
		input_register_b1		: STRING;
		input_register_a0		: STRING;
		multiplier1_direction		: STRING;
		signed_pipeline_aclr_a		: STRING
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (2*mpr-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (2*twr-1 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (twr+mpr DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(twr+mpr DOWNTO 0);
	sub_wire1    <= dataa_0(mpr-1 DOWNTO 0);
	sub_wire3    <= dataa_1(mpr-1 DOWNTO 0);
	sub_wire2    <= sub_wire3(mpr-1 DOWNTO 0) & sub_wire1(mpr-1 DOWNTO 0);
	sub_wire4    <= datab_0(twr-1 DOWNTO 0);
	sub_wire6    <= datab_1(twr-1 DOWNTO 0);
	sub_wire5    <= sub_wire6(twr-1 DOWNTO 0) & sub_wire4(twr-1 DOWNTO 0);

	ALTMULT_ADD_component : altmult_add
	GENERIC MAP (
		input_register_a1 => "CLOCK0",
		multiplier_register0 => "CLOCK0",
		signed_pipeline_aclr_b => "UNUSED",
		multiplier_register1 => "CLOCK0",
		addnsub_multiplier_pipeline_aclr1 => "UNUSED",
		signed_aclr_a => "UNUSED",
		signed_register_a => "CLOCK0",
		number_of_multipliers => 2,
		multiplier_aclr0 => "UNUSED",
		signed_aclr_b => "UNUSED",
		signed_register_b => "CLOCK0",
		lpm_type => "altmult_add",
		multiplier_aclr1 => "UNUSED",
		input_aclr_b0 => "UNUSED",
		output_register => "CLOCK0",
		representation_a => "SIGNED",
		signed_pipeline_register_a => "CLOCK0",
		width_result => mpr+twr+1,
		input_source_b0 => "DATAB",
		input_aclr_b1 => "UNUSED",
		input_aclr_a0 => "UNUSED",
		addnsub_multiplier_register1 => "CLOCK0",
		representation_b => "SIGNED",
		signed_pipeline_register_b => "CLOCK0",
		input_source_b1 => "DATAB",
		input_source_a0 => "DATAA",
		input_aclr_a1 => "UNUSED",
		dedicated_multiplier_circuitry => "AUTO",
		input_source_a1 => "DATAA",
		addnsub_multiplier_aclr1 => "UNUSED",
		output_aclr => "UNUSED",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		width_a => mpr,
		input_register_b0 => "CLOCK0",
		width_b => twr,
		input_register_b1 => "CLOCK0",
		input_register_a0 => "CLOCK0",
		multiplier1_direction => dirn,
		signed_pipeline_aclr_a => "UNUSED"
	)
	PORT MAP (
		dataa => sub_wire2,
		datab => sub_wire5,
		clock0 => clock0,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: SRCA0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNA STRING "Signed"
-- Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: MULT_REGOUT0 STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB STRING "Signed"
-- Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: SAME_CONFIG STRING "1"
-- Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGB0 STRING "1"
-- Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGA0 STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED STRING "0"
-- Retrieval info: PRIVATE: RTS_WIDTH STRING "29"
-- Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: IMPL_STYLE_LCELL STRING "0"
-- Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: NUM_MULT STRING "2"
-- Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: SCANOUTA STRING "0"
-- Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: REG_OUT STRING "1"
-- Retrieval info: PRIVATE: SCANOUTB STRING "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT STRING "1"
-- Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADD_ENABLE STRING "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ALL_REG_ACLR STRING "0"
-- Retrieval info: PRIVATE: WIDTHA STRING "16"
-- Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_REG STRING "1"
-- Retrieval info: PRIVATE: WIDTHB STRING "12"
-- Retrieval info: PRIVATE: SIGNB_REG STRING "1"
-- Retrieval info: PRIVATE: OP1 STRING "Subtract"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB1_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: OP3 STRING "Add"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INPUT_REGISTER_A1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_B STRING "UNUSED"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_ACLR1 STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGNED_ACLR_A STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: NUMBER_OF_MULTIPLIERS NUMERIC "2"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR0 STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGNED_ACLR_B STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_add"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR1 STRING "UNUSED"
-- Retrieval info: CONSTANT: INPUT_ACLR_B0 STRING "UNUSED"
-- Retrieval info: CONSTANT: OUTPUT_REGISTER STRING "CLOCK0"
-- Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "29"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B0 STRING "DATAB"
-- Retrieval info: CONSTANT: INPUT_ACLR_B1 STRING "UNUSED"
-- Retrieval info: CONSTANT: INPUT_ACLR_A0 STRING "UNUSED"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B1 STRING "DATAB"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A0 STRING "DATAA"
-- Retrieval info: CONSTANT: INPUT_ACLR_A1 STRING "UNUSED"
-- Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "AUTO"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A1 STRING "DATAA"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_ACLR1 STRING "UNUSED"
-- Retrieval info: CONSTANT: OUTPUT_ACLR STRING "UNUSED"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "12"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER1_DIRECTION STRING "SUB"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_A STRING "UNUSED"
-- Retrieval info: USED_PORT: clock0 0 0 0 0 INPUT VCC "clock0"
-- Retrieval info: USED_PORT: dataa_0 0 0 16 0 INPUT GND "dataa_0[15..0]"
-- Retrieval info: USED_PORT: dataa_1 0 0 16 0 INPUT GND "dataa_1[15..0]"
-- Retrieval info: USED_PORT: datab_0 0 0 12 0 INPUT GND "datab_0[11..0]"
-- Retrieval info: USED_PORT: datab_1 0 0 12 0 INPUT GND "datab_1[11..0]"
-- Retrieval info: USED_PORT: result 0 0 29 0 OUTPUT GND "result[28..0]"
-- Retrieval info: CONNECT: @datab 0 0 12 12 datab_1 0 0 12 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock0 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 29 0 @result 0 0 29 0
-- Retrieval info: CONNECT: @dataa 0 0 16 0 dataa_0 0 0 16 0
-- Retrieval info: CONNECT: @dataa 0 0 16 16 dataa_1 0 0 16 0
-- Retrieval info: CONNECT: @datab 0 0 12 0 datab_0 0 0 12 0
